------------------------------------------------------------------------------
--  Copyright (c) 2018 by Paul Scherrer Institute, Switzerland
--  All rights reserved.
------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

use work.psi_fix_pkg.all;
use work.psi_common_math_pkg.all;

entity psi_fix_lin_approx_inv18b is
  port(
    clk_i : in  std_logic;                         -- system clock
    rst_i : in  std_logic;                         -- system reset
    dat_i : in  std_logic_vector(19 - 1 downto 0); -- Format (0, 1, 18)
    vld_i : in  std_logic;                         -- valid input
    dat_o : out std_logic_vector(18 - 1 downto 0); -- Format (0, 0, 18)
    vld_o : out std_logic                          -- valid output
  );
end entity;

architecture rtl of psi_fix_lin_approx_inv18b is

  -- Constants
  constant InFmt_c      : psi_fix_fmt_t := (0, 1, 18);
  constant OutFmt_c     : psi_fix_fmt_t := (0, 0, 18);
  constant OffsFmt_c    : psi_fix_fmt_t := (1, 0, 21);
  constant GradFmt_c    : psi_fix_fmt_t := (1, 0, 14);
  constant TableSize_c  : integer       := 1024;
  constant TableWidth_c : integer       := 37;

  -- Table

  type Table_t is array (0 to TableSize_c - 1) of std_logic_vector(TableWidth_c - 1 downto 0);
  constant Table_c : Table_t := (
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16384, 15) & to_signed(2097151, 22)),
    std_logic_vector(to_signed(-16352, 15) & to_signed(2095106, 22)),
    std_logic_vector(to_signed(-16288, 15) & to_signed(2091026, 22)),
    std_logic_vector(to_signed(-16225, 15) & to_signed(2086962, 22)),
    std_logic_vector(to_signed(-16162, 15) & to_signed(2082913, 22)),
    std_logic_vector(to_signed(-16100, 15) & to_signed(2078881, 22)),
    std_logic_vector(to_signed(-16038, 15) & to_signed(2074863, 22)),
    std_logic_vector(to_signed(-15976, 15) & to_signed(2070862, 22)),
    std_logic_vector(to_signed(-15914, 15) & to_signed(2066876, 22)),
    std_logic_vector(to_signed(-15853, 15) & to_signed(2062905, 22)),
    std_logic_vector(to_signed(-15793, 15) & to_signed(2058949, 22)),
    std_logic_vector(to_signed(-15732, 15) & to_signed(2055008, 22)),
    std_logic_vector(to_signed(-15672, 15) & to_signed(2051083, 22)),
    std_logic_vector(to_signed(-15612, 15) & to_signed(2047172, 22)),
    std_logic_vector(to_signed(-15553, 15) & to_signed(2043277, 22)),
    std_logic_vector(to_signed(-15494, 15) & to_signed(2039396, 22)),
    std_logic_vector(to_signed(-15435, 15) & to_signed(2035530, 22)),
    std_logic_vector(to_signed(-15377, 15) & to_signed(2031678, 22)),
    std_logic_vector(to_signed(-15319, 15) & to_signed(2027841, 22)),
    std_logic_vector(to_signed(-15261, 15) & to_signed(2024019, 22)),
    std_logic_vector(to_signed(-15204, 15) & to_signed(2020210, 22)),
    std_logic_vector(to_signed(-15147, 15) & to_signed(2016417, 22)),
    std_logic_vector(to_signed(-15090, 15) & to_signed(2012637, 22)),
    std_logic_vector(to_signed(-15034, 15) & to_signed(2008872, 22)),
    std_logic_vector(to_signed(-14978, 15) & to_signed(2005120, 22)),
    std_logic_vector(to_signed(-14922, 15) & to_signed(2001383, 22)),
    std_logic_vector(to_signed(-14866, 15) & to_signed(1997659, 22)),
    std_logic_vector(to_signed(-14811, 15) & to_signed(1993950, 22)),
    std_logic_vector(to_signed(-14756, 15) & to_signed(1990254, 22)),
    std_logic_vector(to_signed(-14702, 15) & to_signed(1986571, 22)),
    std_logic_vector(to_signed(-14647, 15) & to_signed(1982903, 22)),
    std_logic_vector(to_signed(-14594, 15) & to_signed(1979248, 22)),
    std_logic_vector(to_signed(-14540, 15) & to_signed(1975606, 22)),
    std_logic_vector(to_signed(-14487, 15) & to_signed(1971978, 22)),
    std_logic_vector(to_signed(-14433, 15) & to_signed(1968363, 22)),
    std_logic_vector(to_signed(-14381, 15) & to_signed(1964761, 22)),
    std_logic_vector(to_signed(-14328, 15) & to_signed(1961172, 22)),
    std_logic_vector(to_signed(-14276, 15) & to_signed(1957597, 22)),
    std_logic_vector(to_signed(-14224, 15) & to_signed(1954034, 22)),
    std_logic_vector(to_signed(-14172, 15) & to_signed(1950485, 22)),
    std_logic_vector(to_signed(-14121, 15) & to_signed(1946948, 22)),
    std_logic_vector(to_signed(-14070, 15) & to_signed(1943424, 22)),
    std_logic_vector(to_signed(-14019, 15) & to_signed(1939913, 22)),
    std_logic_vector(to_signed(-13969, 15) & to_signed(1936414, 22)),
    std_logic_vector(to_signed(-13918, 15) & to_signed(1932929, 22)),
    std_logic_vector(to_signed(-13869, 15) & to_signed(1929455, 22)),
    std_logic_vector(to_signed(-13819, 15) & to_signed(1925994, 22)),
    std_logic_vector(to_signed(-13769, 15) & to_signed(1922546, 22)),
    std_logic_vector(to_signed(-13720, 15) & to_signed(1919110, 22)),
    std_logic_vector(to_signed(-13671, 15) & to_signed(1915686, 22)),
    std_logic_vector(to_signed(-13623, 15) & to_signed(1912274, 22)),
    std_logic_vector(to_signed(-13574, 15) & to_signed(1908874, 22)),
    std_logic_vector(to_signed(-13526, 15) & to_signed(1905487, 22)),
    std_logic_vector(to_signed(-13478, 15) & to_signed(1902111, 22)),
    std_logic_vector(to_signed(-13431, 15) & to_signed(1898748, 22)),
    std_logic_vector(to_signed(-13383, 15) & to_signed(1895396, 22)),
    std_logic_vector(to_signed(-13336, 15) & to_signed(1892056, 22)),
    std_logic_vector(to_signed(-13289, 15) & to_signed(1888728, 22)),
    std_logic_vector(to_signed(-13243, 15) & to_signed(1885411, 22)),
    std_logic_vector(to_signed(-13196, 15) & to_signed(1882107, 22)),
    std_logic_vector(to_signed(-13150, 15) & to_signed(1878813, 22)),
    std_logic_vector(to_signed(-13104, 15) & to_signed(1875532, 22)),
    std_logic_vector(to_signed(-13058, 15) & to_signed(1872261, 22)),
    std_logic_vector(to_signed(-13013, 15) & to_signed(1869002, 22)),
    std_logic_vector(to_signed(-12968, 15) & to_signed(1865755, 22)),
    std_logic_vector(to_signed(-12923, 15) & to_signed(1862518, 22)),
    std_logic_vector(to_signed(-12878, 15) & to_signed(1859293, 22)),
    std_logic_vector(to_signed(-12834, 15) & to_signed(1856079, 22)),
    std_logic_vector(to_signed(-12789, 15) & to_signed(1852876, 22)),
    std_logic_vector(to_signed(-12745, 15) & to_signed(1849684, 22)),
    std_logic_vector(to_signed(-12702, 15) & to_signed(1846504, 22)),
    std_logic_vector(to_signed(-12658, 15) & to_signed(1843334, 22)),
    std_logic_vector(to_signed(-12615, 15) & to_signed(1840175, 22)),
    std_logic_vector(to_signed(-12572, 15) & to_signed(1837026, 22)),
    std_logic_vector(to_signed(-12529, 15) & to_signed(1833889, 22)),
    std_logic_vector(to_signed(-12486, 15) & to_signed(1830762, 22)),
    std_logic_vector(to_signed(-12444, 15) & to_signed(1827646, 22)),
    std_logic_vector(to_signed(-12401, 15) & to_signed(1824540, 22)),
    std_logic_vector(to_signed(-12359, 15) & to_signed(1821445, 22)),
    std_logic_vector(to_signed(-12317, 15) & to_signed(1818360, 22)),
    std_logic_vector(to_signed(-12276, 15) & to_signed(1815286, 22)),
    std_logic_vector(to_signed(-12234, 15) & to_signed(1812222, 22)),
    std_logic_vector(to_signed(-12193, 15) & to_signed(1809169, 22)),
    std_logic_vector(to_signed(-12152, 15) & to_signed(1806126, 22)),
    std_logic_vector(to_signed(-12111, 15) & to_signed(1803093, 22)),
    std_logic_vector(to_signed(-12071, 15) & to_signed(1800070, 22)),
    std_logic_vector(to_signed(-12031, 15) & to_signed(1797057, 22)),
    std_logic_vector(to_signed(-11990, 15) & to_signed(1794055, 22)),
    std_logic_vector(to_signed(-11950, 15) & to_signed(1791062, 22)),
    std_logic_vector(to_signed(-11911, 15) & to_signed(1788080, 22)),
    std_logic_vector(to_signed(-11871, 15) & to_signed(1785107, 22)),
    std_logic_vector(to_signed(-11832, 15) & to_signed(1782144, 22)),
    std_logic_vector(to_signed(-11792, 15) & to_signed(1779191, 22)),
    std_logic_vector(to_signed(-11754, 15) & to_signed(1776248, 22)),
    std_logic_vector(to_signed(-11715, 15) & to_signed(1773314, 22)),
    std_logic_vector(to_signed(-11676, 15) & to_signed(1770390, 22)),
    std_logic_vector(to_signed(-11638, 15) & to_signed(1767476, 22)),
    std_logic_vector(to_signed(-11599, 15) & to_signed(1764572, 22)),
    std_logic_vector(to_signed(-11561, 15) & to_signed(1761676, 22)),
    std_logic_vector(to_signed(-11524, 15) & to_signed(1758791, 22)),
    std_logic_vector(to_signed(-11486, 15) & to_signed(1755915, 22)),
    std_logic_vector(to_signed(-11448, 15) & to_signed(1753048, 22)),
    std_logic_vector(to_signed(-11411, 15) & to_signed(1750190, 22)),
    std_logic_vector(to_signed(-11374, 15) & to_signed(1747342, 22)),
    std_logic_vector(to_signed(-11337, 15) & to_signed(1744503, 22)),
    std_logic_vector(to_signed(-11300, 15) & to_signed(1741674, 22)),
    std_logic_vector(to_signed(-11264, 15) & to_signed(1738853, 22)),
    std_logic_vector(to_signed(-11227, 15) & to_signed(1736042, 22)),
    std_logic_vector(to_signed(-11191, 15) & to_signed(1733239, 22)),
    std_logic_vector(to_signed(-11155, 15) & to_signed(1730446, 22)),
    std_logic_vector(to_signed(-11119, 15) & to_signed(1727662, 22)),
    std_logic_vector(to_signed(-11084, 15) & to_signed(1724886, 22)),
    std_logic_vector(to_signed(-11048, 15) & to_signed(1722120, 22)),
    std_logic_vector(to_signed(-11013, 15) & to_signed(1719362, 22)),
    std_logic_vector(to_signed(-10978, 15) & to_signed(1716614, 22)),
    std_logic_vector(to_signed(-10943, 15) & to_signed(1713874, 22)),
    std_logic_vector(to_signed(-10908, 15) & to_signed(1711142, 22)),
    std_logic_vector(to_signed(-10873, 15) & to_signed(1708420, 22)),
    std_logic_vector(to_signed(-10838, 15) & to_signed(1705706, 22)),
    std_logic_vector(to_signed(-10804, 15) & to_signed(1703001, 22)),
    std_logic_vector(to_signed(-10770, 15) & to_signed(1700304, 22)),
    std_logic_vector(to_signed(-10736, 15) & to_signed(1697616, 22)),
    std_logic_vector(to_signed(-10702, 15) & to_signed(1694936, 22)),
    std_logic_vector(to_signed(-10668, 15) & to_signed(1692264, 22)),
    std_logic_vector(to_signed(-10635, 15) & to_signed(1689602, 22)),
    std_logic_vector(to_signed(-10601, 15) & to_signed(1686947, 22)),
    std_logic_vector(to_signed(-10568, 15) & to_signed(1684301, 22)),
    std_logic_vector(to_signed(-10535, 15) & to_signed(1681663, 22)),
    std_logic_vector(to_signed(-10502, 15) & to_signed(1679033, 22)),
    std_logic_vector(to_signed(-10469, 15) & to_signed(1676412, 22)),
    std_logic_vector(to_signed(-10437, 15) & to_signed(1673799, 22)),
    std_logic_vector(to_signed(-10404, 15) & to_signed(1671194, 22)),
    std_logic_vector(to_signed(-10372, 15) & to_signed(1668596, 22)),
    std_logic_vector(to_signed(-10340, 15) & to_signed(1666007, 22)),
    std_logic_vector(to_signed(-10308, 15) & to_signed(1663427, 22)),
    std_logic_vector(to_signed(-10276, 15) & to_signed(1660854, 22)),
    std_logic_vector(to_signed(-10244, 15) & to_signed(1658289, 22)),
    std_logic_vector(to_signed(-10213, 15) & to_signed(1655731, 22)),
    std_logic_vector(to_signed(-10181, 15) & to_signed(1653182, 22)),
    std_logic_vector(to_signed(-10150, 15) & to_signed(1650641, 22)),
    std_logic_vector(to_signed(-10119, 15) & to_signed(1648107, 22)),
    std_logic_vector(to_signed(-10088, 15) & to_signed(1645581, 22)),
    std_logic_vector(to_signed(-10057, 15) & to_signed(1643063, 22)),
    std_logic_vector(to_signed(-10026, 15) & to_signed(1640553, 22)),
    std_logic_vector(to_signed(-9996, 15) & to_signed(1638050, 22)),
    std_logic_vector(to_signed(-9965, 15) & to_signed(1635555, 22)),
    std_logic_vector(to_signed(-9935, 15) & to_signed(1633067, 22)),
    std_logic_vector(to_signed(-9905, 15) & to_signed(1630587, 22)),
    std_logic_vector(to_signed(-9875, 15) & to_signed(1628115, 22)),
    std_logic_vector(to_signed(-9845, 15) & to_signed(1625650, 22)),
    std_logic_vector(to_signed(-9815, 15) & to_signed(1623192, 22)),
    std_logic_vector(to_signed(-9786, 15) & to_signed(1620742, 22)),
    std_logic_vector(to_signed(-9756, 15) & to_signed(1618300, 22)),
    std_logic_vector(to_signed(-9727, 15) & to_signed(1615864, 22)),
    std_logic_vector(to_signed(-9698, 15) & to_signed(1613436, 22)),
    std_logic_vector(to_signed(-9669, 15) & to_signed(1611015, 22)),
    std_logic_vector(to_signed(-9640, 15) & to_signed(1608602, 22)),
    std_logic_vector(to_signed(-9611, 15) & to_signed(1606196, 22)),
    std_logic_vector(to_signed(-9582, 15) & to_signed(1603797, 22)),
    std_logic_vector(to_signed(-9553, 15) & to_signed(1601405, 22)),
    std_logic_vector(to_signed(-9525, 15) & to_signed(1599020, 22)),
    std_logic_vector(to_signed(-9497, 15) & to_signed(1596642, 22)),
    std_logic_vector(to_signed(-9469, 15) & to_signed(1594271, 22)),
    std_logic_vector(to_signed(-9441, 15) & to_signed(1591908, 22)),
    std_logic_vector(to_signed(-9413, 15) & to_signed(1589551, 22)),
    std_logic_vector(to_signed(-9385, 15) & to_signed(1587202, 22)),
    std_logic_vector(to_signed(-9357, 15) & to_signed(1584859, 22)),
    std_logic_vector(to_signed(-9330, 15) & to_signed(1582523, 22)),
    std_logic_vector(to_signed(-9302, 15) & to_signed(1580194, 22)),
    std_logic_vector(to_signed(-9275, 15) & to_signed(1577872, 22)),
    std_logic_vector(to_signed(-9248, 15) & to_signed(1575557, 22)),
    std_logic_vector(to_signed(-9221, 15) & to_signed(1573248, 22)),
    std_logic_vector(to_signed(-9194, 15) & to_signed(1570946, 22)),
    std_logic_vector(to_signed(-9167, 15) & to_signed(1568651, 22)),
    std_logic_vector(to_signed(-9140, 15) & to_signed(1566363, 22)),
    std_logic_vector(to_signed(-9113, 15) & to_signed(1564081, 22)),
    std_logic_vector(to_signed(-9087, 15) & to_signed(1561806, 22)),
    std_logic_vector(to_signed(-9060, 15) & to_signed(1559538, 22)),
    std_logic_vector(to_signed(-9034, 15) & to_signed(1557276, 22)),
    std_logic_vector(to_signed(-9008, 15) & to_signed(1555021, 22)),
    std_logic_vector(to_signed(-8982, 15) & to_signed(1552772, 22)),
    std_logic_vector(to_signed(-8956, 15) & to_signed(1550530, 22)),
    std_logic_vector(to_signed(-8930, 15) & to_signed(1548294, 22)),
    std_logic_vector(to_signed(-8905, 15) & to_signed(1546065, 22)),
    std_logic_vector(to_signed(-8879, 15) & to_signed(1543842, 22)),
    std_logic_vector(to_signed(-8854, 15) & to_signed(1541625, 22)),
    std_logic_vector(to_signed(-8828, 15) & to_signed(1539415, 22)),
    std_logic_vector(to_signed(-8803, 15) & to_signed(1537211, 22)),
    std_logic_vector(to_signed(-8778, 15) & to_signed(1535013, 22)),
    std_logic_vector(to_signed(-8753, 15) & to_signed(1532822, 22)),
    std_logic_vector(to_signed(-8728, 15) & to_signed(1530637, 22)),
    std_logic_vector(to_signed(-8703, 15) & to_signed(1528458, 22)),
    std_logic_vector(to_signed(-8678, 15) & to_signed(1526285, 22)),
    std_logic_vector(to_signed(-8654, 15) & to_signed(1524119, 22)),
    std_logic_vector(to_signed(-8629, 15) & to_signed(1521959, 22)),
    std_logic_vector(to_signed(-8605, 15) & to_signed(1519804, 22)),
    std_logic_vector(to_signed(-8580, 15) & to_signed(1517656, 22)),
    std_logic_vector(to_signed(-8556, 15) & to_signed(1515514, 22)),
    std_logic_vector(to_signed(-8532, 15) & to_signed(1513378, 22)),
    std_logic_vector(to_signed(-8508, 15) & to_signed(1511248, 22)),
    std_logic_vector(to_signed(-8484, 15) & to_signed(1509124, 22)),
    std_logic_vector(to_signed(-8460, 15) & to_signed(1507006, 22)),
    std_logic_vector(to_signed(-8437, 15) & to_signed(1504894, 22)),
    std_logic_vector(to_signed(-8413, 15) & to_signed(1502788, 22)),
    std_logic_vector(to_signed(-8390, 15) & to_signed(1500687, 22)),
    std_logic_vector(to_signed(-8366, 15) & to_signed(1498593, 22)),
    std_logic_vector(to_signed(-8343, 15) & to_signed(1496504, 22)),
    std_logic_vector(to_signed(-8320, 15) & to_signed(1494421, 22)),
    std_logic_vector(to_signed(-8297, 15) & to_signed(1492344, 22)),
    std_logic_vector(to_signed(-8274, 15) & to_signed(1490273, 22)),
    std_logic_vector(to_signed(-8251, 15) & to_signed(1488208, 22)),
    std_logic_vector(to_signed(-8228, 15) & to_signed(1486148, 22)),
    std_logic_vector(to_signed(-8205, 15) & to_signed(1484094, 22)),
    std_logic_vector(to_signed(-8182, 15) & to_signed(1482045, 22)),
    std_logic_vector(to_signed(-8160, 15) & to_signed(1480003, 22)),
    std_logic_vector(to_signed(-8137, 15) & to_signed(1477965, 22)),
    std_logic_vector(to_signed(-8115, 15) & to_signed(1475934, 22)),
    std_logic_vector(to_signed(-8093, 15) & to_signed(1473908, 22)),
    std_logic_vector(to_signed(-8071, 15) & to_signed(1471887, 22)),
    std_logic_vector(to_signed(-8049, 15) & to_signed(1469872, 22)),
    std_logic_vector(to_signed(-8027, 15) & to_signed(1467863, 22)),
    std_logic_vector(to_signed(-8005, 15) & to_signed(1465859, 22)),
    std_logic_vector(to_signed(-7983, 15) & to_signed(1463861, 22)),
    std_logic_vector(to_signed(-7961, 15) & to_signed(1461868, 22)),
    std_logic_vector(to_signed(-7940, 15) & to_signed(1459880, 22)),
    std_logic_vector(to_signed(-7918, 15) & to_signed(1457898, 22)),
    std_logic_vector(to_signed(-7897, 15) & to_signed(1455921, 22)),
    std_logic_vector(to_signed(-7875, 15) & to_signed(1453950, 22)),
    std_logic_vector(to_signed(-7854, 15) & to_signed(1451984, 22)),
    std_logic_vector(to_signed(-7833, 15) & to_signed(1450023, 22)),
    std_logic_vector(to_signed(-7812, 15) & to_signed(1448067, 22)),
    std_logic_vector(to_signed(-7791, 15) & to_signed(1446117, 22)),
    std_logic_vector(to_signed(-7770, 15) & to_signed(1444172, 22)),
    std_logic_vector(to_signed(-7749, 15) & to_signed(1442232, 22)),
    std_logic_vector(to_signed(-7728, 15) & to_signed(1440298, 22)),
    std_logic_vector(to_signed(-7707, 15) & to_signed(1438368, 22)),
    std_logic_vector(to_signed(-7687, 15) & to_signed(1436444, 22)),
    std_logic_vector(to_signed(-7666, 15) & to_signed(1434525, 22)),
    std_logic_vector(to_signed(-7646, 15) & to_signed(1432611, 22)),
    std_logic_vector(to_signed(-7625, 15) & to_signed(1430702, 22)),
    std_logic_vector(to_signed(-7605, 15) & to_signed(1428798, 22)),
    std_logic_vector(to_signed(-7585, 15) & to_signed(1426899, 22)),
    std_logic_vector(to_signed(-7565, 15) & to_signed(1425006, 22)),
    std_logic_vector(to_signed(-7545, 15) & to_signed(1423117, 22)),
    std_logic_vector(to_signed(-7525, 15) & to_signed(1421233, 22)),
    std_logic_vector(to_signed(-7505, 15) & to_signed(1419355, 22)),
    std_logic_vector(to_signed(-7485, 15) & to_signed(1417481, 22)),
    std_logic_vector(to_signed(-7465, 15) & to_signed(1415612, 22)),
    std_logic_vector(to_signed(-7446, 15) & to_signed(1413748, 22)),
    std_logic_vector(to_signed(-7426, 15) & to_signed(1411889, 22)),
    std_logic_vector(to_signed(-7407, 15) & to_signed(1410035, 22)),
    std_logic_vector(to_signed(-7387, 15) & to_signed(1408186, 22)),
    std_logic_vector(to_signed(-7368, 15) & to_signed(1406342, 22)),
    std_logic_vector(to_signed(-7349, 15) & to_signed(1404502, 22)),
    std_logic_vector(to_signed(-7329, 15) & to_signed(1402667, 22)),
    std_logic_vector(to_signed(-7310, 15) & to_signed(1400837, 22)),
    std_logic_vector(to_signed(-7291, 15) & to_signed(1399012, 22)),
    std_logic_vector(to_signed(-7272, 15) & to_signed(1397192, 22)),
    std_logic_vector(to_signed(-7253, 15) & to_signed(1395376, 22)),
    std_logic_vector(to_signed(-7235, 15) & to_signed(1393565, 22)),
    std_logic_vector(to_signed(-7216, 15) & to_signed(1391759, 22)),
    std_logic_vector(to_signed(-7197, 15) & to_signed(1389957, 22)),
    std_logic_vector(to_signed(-7179, 15) & to_signed(1388160, 22)),
    std_logic_vector(to_signed(-7160, 15) & to_signed(1386368, 22)),
    std_logic_vector(to_signed(-7142, 15) & to_signed(1384580, 22)),
    std_logic_vector(to_signed(-7123, 15) & to_signed(1382797, 22)),
    std_logic_vector(to_signed(-7105, 15) & to_signed(1381018, 22)),
    std_logic_vector(to_signed(-7087, 15) & to_signed(1379244, 22)),
    std_logic_vector(to_signed(-7069, 15) & to_signed(1377475, 22)),
    std_logic_vector(to_signed(-7050, 15) & to_signed(1375710, 22)),
    std_logic_vector(to_signed(-7032, 15) & to_signed(1373950, 22)),
    std_logic_vector(to_signed(-7014, 15) & to_signed(1372194, 22)),
    std_logic_vector(to_signed(-6997, 15) & to_signed(1370443, 22)),
    std_logic_vector(to_signed(-6979, 15) & to_signed(1368696, 22)),
    std_logic_vector(to_signed(-6961, 15) & to_signed(1366953, 22)),
    std_logic_vector(to_signed(-6943, 15) & to_signed(1365215, 22)),
    std_logic_vector(to_signed(-6926, 15) & to_signed(1363482, 22)),
    std_logic_vector(to_signed(-6908, 15) & to_signed(1361752, 22)),
    std_logic_vector(to_signed(-6891, 15) & to_signed(1360028, 22)),
    std_logic_vector(to_signed(-6873, 15) & to_signed(1358307, 22)),
    std_logic_vector(to_signed(-6856, 15) & to_signed(1356591, 22)),
    std_logic_vector(to_signed(-6839, 15) & to_signed(1354879, 22)),
    std_logic_vector(to_signed(-6821, 15) & to_signed(1353172, 22)),
    std_logic_vector(to_signed(-6804, 15) & to_signed(1351469, 22)),
    std_logic_vector(to_signed(-6787, 15) & to_signed(1349770, 22)),
    std_logic_vector(to_signed(-6770, 15) & to_signed(1348075, 22)),
    std_logic_vector(to_signed(-6753, 15) & to_signed(1346385, 22)),
    std_logic_vector(to_signed(-6736, 15) & to_signed(1344699, 22)),
    std_logic_vector(to_signed(-6719, 15) & to_signed(1343017, 22)),
    std_logic_vector(to_signed(-6703, 15) & to_signed(1341339, 22)),
    std_logic_vector(to_signed(-6686, 15) & to_signed(1339665, 22)),
    std_logic_vector(to_signed(-6669, 15) & to_signed(1337996, 22)),
    std_logic_vector(to_signed(-6653, 15) & to_signed(1336331, 22)),
    std_logic_vector(to_signed(-6636, 15) & to_signed(1334670, 22)),
    std_logic_vector(to_signed(-6620, 15) & to_signed(1333013, 22)),
    std_logic_vector(to_signed(-6603, 15) & to_signed(1331360, 22)),
    std_logic_vector(to_signed(-6587, 15) & to_signed(1329711, 22)),
    std_logic_vector(to_signed(-6571, 15) & to_signed(1328067, 22)),
    std_logic_vector(to_signed(-6554, 15) & to_signed(1326426, 22)),
    std_logic_vector(to_signed(-6538, 15) & to_signed(1324789, 22)),
    std_logic_vector(to_signed(-6522, 15) & to_signed(1323157, 22)),
    std_logic_vector(to_signed(-6506, 15) & to_signed(1321528, 22)),
    std_logic_vector(to_signed(-6490, 15) & to_signed(1319904, 22)),
    std_logic_vector(to_signed(-6474, 15) & to_signed(1318283, 22)),
    std_logic_vector(to_signed(-6458, 15) & to_signed(1316667, 22)),
    std_logic_vector(to_signed(-6442, 15) & to_signed(1315054, 22)),
    std_logic_vector(to_signed(-6427, 15) & to_signed(1313446, 22)),
    std_logic_vector(to_signed(-6411, 15) & to_signed(1311841, 22)),
    std_logic_vector(to_signed(-6395, 15) & to_signed(1310240, 22)),
    std_logic_vector(to_signed(-6380, 15) & to_signed(1308643, 22)),
    std_logic_vector(to_signed(-6364, 15) & to_signed(1307050, 22)),
    std_logic_vector(to_signed(-6349, 15) & to_signed(1305461, 22)),
    std_logic_vector(to_signed(-6333, 15) & to_signed(1303876, 22)),
    std_logic_vector(to_signed(-6318, 15) & to_signed(1302295, 22)),
    std_logic_vector(to_signed(-6303, 15) & to_signed(1300717, 22)),
    std_logic_vector(to_signed(-6287, 15) & to_signed(1299143, 22)),
    std_logic_vector(to_signed(-6272, 15) & to_signed(1297573, 22)),
    std_logic_vector(to_signed(-6257, 15) & to_signed(1296007, 22)),
    std_logic_vector(to_signed(-6242, 15) & to_signed(1294445, 22)),
    std_logic_vector(to_signed(-6227, 15) & to_signed(1292886, 22)),
    std_logic_vector(to_signed(-6212, 15) & to_signed(1291331, 22)),
    std_logic_vector(to_signed(-6197, 15) & to_signed(1289780, 22)),
    std_logic_vector(to_signed(-6182, 15) & to_signed(1288233, 22)),
    std_logic_vector(to_signed(-6167, 15) & to_signed(1286689, 22)),
    std_logic_vector(to_signed(-6153, 15) & to_signed(1285149, 22)),
    std_logic_vector(to_signed(-6138, 15) & to_signed(1283612, 22)),
    std_logic_vector(to_signed(-6123, 15) & to_signed(1282080, 22)),
    std_logic_vector(to_signed(-6109, 15) & to_signed(1280551, 22)),
    std_logic_vector(to_signed(-6094, 15) & to_signed(1279025, 22)),
    std_logic_vector(to_signed(-6080, 15) & to_signed(1277504, 22)),
    std_logic_vector(to_signed(-6065, 15) & to_signed(1275986, 22)),
    std_logic_vector(to_signed(-6051, 15) & to_signed(1274471, 22)),
    std_logic_vector(to_signed(-6037, 15) & to_signed(1272960, 22)),
    std_logic_vector(to_signed(-6022, 15) & to_signed(1271453, 22)),
    std_logic_vector(to_signed(-6008, 15) & to_signed(1269949, 22)),
    std_logic_vector(to_signed(-5994, 15) & to_signed(1268449, 22)),
    std_logic_vector(to_signed(-5980, 15) & to_signed(1266952, 22)),
    std_logic_vector(to_signed(-5966, 15) & to_signed(1265459, 22)),
    std_logic_vector(to_signed(-5952, 15) & to_signed(1263969, 22)),
    std_logic_vector(to_signed(-5938, 15) & to_signed(1262483, 22)),
    std_logic_vector(to_signed(-5924, 15) & to_signed(1261000, 22)),
    std_logic_vector(to_signed(-5910, 15) & to_signed(1259521, 22)),
    std_logic_vector(to_signed(-5896, 15) & to_signed(1258045, 22)),
    std_logic_vector(to_signed(-5882, 15) & to_signed(1256573, 22)),
    std_logic_vector(to_signed(-5868, 15) & to_signed(1255104, 22)),
    std_logic_vector(to_signed(-5855, 15) & to_signed(1253639, 22)),
    std_logic_vector(to_signed(-5841, 15) & to_signed(1252177, 22)),
    std_logic_vector(to_signed(-5827, 15) & to_signed(1250718, 22)),
    std_logic_vector(to_signed(-5814, 15) & to_signed(1249263, 22)),
    std_logic_vector(to_signed(-5800, 15) & to_signed(1247812, 22)),
    std_logic_vector(to_signed(-5787, 15) & to_signed(1246363, 22)),
    std_logic_vector(to_signed(-5774, 15) & to_signed(1244918, 22)),
    std_logic_vector(to_signed(-5760, 15) & to_signed(1243476, 22)),
    std_logic_vector(to_signed(-5747, 15) & to_signed(1242038, 22)),
    std_logic_vector(to_signed(-5734, 15) & to_signed(1240603, 22)),
    std_logic_vector(to_signed(-5720, 15) & to_signed(1239171, 22)),
    std_logic_vector(to_signed(-5707, 15) & to_signed(1237743, 22)),
    std_logic_vector(to_signed(-5694, 15) & to_signed(1236318, 22)),
    std_logic_vector(to_signed(-5681, 15) & to_signed(1234896, 22)),
    std_logic_vector(to_signed(-5668, 15) & to_signed(1233477, 22)),
    std_logic_vector(to_signed(-5655, 15) & to_signed(1232062, 22)),
    std_logic_vector(to_signed(-5642, 15) & to_signed(1230650, 22)),
    std_logic_vector(to_signed(-5629, 15) & to_signed(1229241, 22)),
    std_logic_vector(to_signed(-5616, 15) & to_signed(1227835, 22)),
    std_logic_vector(to_signed(-5603, 15) & to_signed(1226433, 22)),
    std_logic_vector(to_signed(-5591, 15) & to_signed(1225033, 22)),
    std_logic_vector(to_signed(-5578, 15) & to_signed(1223637, 22)),
    std_logic_vector(to_signed(-5565, 15) & to_signed(1222245, 22)),
    std_logic_vector(to_signed(-5552, 15) & to_signed(1220855, 22)),
    std_logic_vector(to_signed(-5540, 15) & to_signed(1219468, 22)),
    std_logic_vector(to_signed(-5527, 15) & to_signed(1218085, 22)),
    std_logic_vector(to_signed(-5515, 15) & to_signed(1216705, 22)),
    std_logic_vector(to_signed(-5502, 15) & to_signed(1215327, 22)),
    std_logic_vector(to_signed(-5490, 15) & to_signed(1213953, 22)),
    std_logic_vector(to_signed(-5478, 15) & to_signed(1212583, 22)),
    std_logic_vector(to_signed(-5465, 15) & to_signed(1211215, 22)),
    std_logic_vector(to_signed(-5453, 15) & to_signed(1209850, 22)),
    std_logic_vector(to_signed(-5441, 15) & to_signed(1208488, 22)),
    std_logic_vector(to_signed(-5428, 15) & to_signed(1207130, 22)),
    std_logic_vector(to_signed(-5416, 15) & to_signed(1205774, 22)),
    std_logic_vector(to_signed(-5404, 15) & to_signed(1204422, 22)),
    std_logic_vector(to_signed(-5392, 15) & to_signed(1203072, 22)),
    std_logic_vector(to_signed(-5380, 15) & to_signed(1201726, 22)),
    std_logic_vector(to_signed(-5368, 15) & to_signed(1200382, 22)),
    std_logic_vector(to_signed(-5356, 15) & to_signed(1199042, 22)),
    std_logic_vector(to_signed(-5344, 15) & to_signed(1197704, 22)),
    std_logic_vector(to_signed(-5332, 15) & to_signed(1196370, 22)),
    std_logic_vector(to_signed(-5320, 15) & to_signed(1195038, 22)),
    std_logic_vector(to_signed(-5308, 15) & to_signed(1193710, 22)),
    std_logic_vector(to_signed(-5297, 15) & to_signed(1192384, 22)),
    std_logic_vector(to_signed(-5285, 15) & to_signed(1191061, 22)),
    std_logic_vector(to_signed(-5273, 15) & to_signed(1189742, 22)),
    std_logic_vector(to_signed(-5261, 15) & to_signed(1188425, 22)),
    std_logic_vector(to_signed(-5250, 15) & to_signed(1187111, 22)),
    std_logic_vector(to_signed(-5238, 15) & to_signed(1185800, 22)),
    std_logic_vector(to_signed(-5227, 15) & to_signed(1184492, 22)),
    std_logic_vector(to_signed(-5215, 15) & to_signed(1183187, 22)),
    std_logic_vector(to_signed(-5204, 15) & to_signed(1181884, 22)),
    std_logic_vector(to_signed(-5192, 15) & to_signed(1180585, 22)),
    std_logic_vector(to_signed(-5181, 15) & to_signed(1179288, 22)),
    std_logic_vector(to_signed(-5169, 15) & to_signed(1177994, 22)),
    std_logic_vector(to_signed(-5158, 15) & to_signed(1176703, 22)),
    std_logic_vector(to_signed(-5147, 15) & to_signed(1175415, 22)),
    std_logic_vector(to_signed(-5136, 15) & to_signed(1174130, 22)),
    std_logic_vector(to_signed(-5124, 15) & to_signed(1172847, 22)),
    std_logic_vector(to_signed(-5113, 15) & to_signed(1171568, 22)),
    std_logic_vector(to_signed(-5102, 15) & to_signed(1170291, 22)),
    std_logic_vector(to_signed(-5091, 15) & to_signed(1169017, 22)),
    std_logic_vector(to_signed(-5080, 15) & to_signed(1167745, 22)),
    std_logic_vector(to_signed(-5069, 15) & to_signed(1166477, 22)),
    std_logic_vector(to_signed(-5058, 15) & to_signed(1165211, 22)),
    std_logic_vector(to_signed(-5047, 15) & to_signed(1163948, 22)),
    std_logic_vector(to_signed(-5036, 15) & to_signed(1162687, 22)),
    std_logic_vector(to_signed(-5025, 15) & to_signed(1161430, 22)),
    std_logic_vector(to_signed(-5014, 15) & to_signed(1160175, 22)),
    std_logic_vector(to_signed(-5003, 15) & to_signed(1158923, 22)),
    std_logic_vector(to_signed(-4993, 15) & to_signed(1157673, 22)),
    std_logic_vector(to_signed(-4982, 15) & to_signed(1156426, 22)),
    std_logic_vector(to_signed(-4971, 15) & to_signed(1155182, 22)),
    std_logic_vector(to_signed(-4961, 15) & to_signed(1153941, 22)),
    std_logic_vector(to_signed(-4950, 15) & to_signed(1152702, 22)),
    std_logic_vector(to_signed(-4939, 15) & to_signed(1151466, 22)),
    std_logic_vector(to_signed(-4929, 15) & to_signed(1150232, 22)),
    std_logic_vector(to_signed(-4918, 15) & to_signed(1149001, 22)),
    std_logic_vector(to_signed(-4908, 15) & to_signed(1147773, 22)),
    std_logic_vector(to_signed(-4897, 15) & to_signed(1146548, 22)),
    std_logic_vector(to_signed(-4887, 15) & to_signed(1145325, 22)),
    std_logic_vector(to_signed(-4876, 15) & to_signed(1144104, 22)),
    std_logic_vector(to_signed(-4866, 15) & to_signed(1142886, 22)),
    std_logic_vector(to_signed(-4856, 15) & to_signed(1141671, 22)),
    std_logic_vector(to_signed(-4845, 15) & to_signed(1140459, 22)),
    std_logic_vector(to_signed(-4835, 15) & to_signed(1139249, 22)),
    std_logic_vector(to_signed(-4825, 15) & to_signed(1138041, 22)),
    std_logic_vector(to_signed(-4815, 15) & to_signed(1136836, 22)),
    std_logic_vector(to_signed(-4804, 15) & to_signed(1135634, 22)),
    std_logic_vector(to_signed(-4794, 15) & to_signed(1134434, 22)),
    std_logic_vector(to_signed(-4784, 15) & to_signed(1133237, 22)),
    std_logic_vector(to_signed(-4774, 15) & to_signed(1132042, 22)),
    std_logic_vector(to_signed(-4764, 15) & to_signed(1130850, 22)),
    std_logic_vector(to_signed(-4754, 15) & to_signed(1129660, 22)),
    std_logic_vector(to_signed(-4744, 15) & to_signed(1128473, 22)),
    std_logic_vector(to_signed(-4734, 15) & to_signed(1127288, 22)),
    std_logic_vector(to_signed(-4724, 15) & to_signed(1126106, 22)),
    std_logic_vector(to_signed(-4714, 15) & to_signed(1124926, 22)),
    std_logic_vector(to_signed(-4704, 15) & to_signed(1123749, 22)),
    std_logic_vector(to_signed(-4695, 15) & to_signed(1122574, 22)),
    std_logic_vector(to_signed(-4685, 15) & to_signed(1121401, 22)),
    std_logic_vector(to_signed(-4675, 15) & to_signed(1120231, 22)),
    std_logic_vector(to_signed(-4665, 15) & to_signed(1119064, 22)),
    std_logic_vector(to_signed(-4655, 15) & to_signed(1117899, 22)),
    std_logic_vector(to_signed(-4646, 15) & to_signed(1116736, 22)),
    std_logic_vector(to_signed(-4636, 15) & to_signed(1115576, 22)),
    std_logic_vector(to_signed(-4627, 15) & to_signed(1114418, 22)),
    std_logic_vector(to_signed(-4617, 15) & to_signed(1113263, 22)),
    std_logic_vector(to_signed(-4607, 15) & to_signed(1112110, 22)),
    std_logic_vector(to_signed(-4598, 15) & to_signed(1110959, 22)),
    std_logic_vector(to_signed(-4588, 15) & to_signed(1109811, 22)),
    std_logic_vector(to_signed(-4579, 15) & to_signed(1108665, 22)),
    std_logic_vector(to_signed(-4569, 15) & to_signed(1107521, 22)),
    std_logic_vector(to_signed(-4560, 15) & to_signed(1106380, 22)),
    std_logic_vector(to_signed(-4551, 15) & to_signed(1105241, 22)),
    std_logic_vector(to_signed(-4541, 15) & to_signed(1104105, 22)),
    std_logic_vector(to_signed(-4532, 15) & to_signed(1102971, 22)),
    std_logic_vector(to_signed(-4523, 15) & to_signed(1101839, 22)),
    std_logic_vector(to_signed(-4513, 15) & to_signed(1100709, 22)),
    std_logic_vector(to_signed(-4504, 15) & to_signed(1099582, 22)),
    std_logic_vector(to_signed(-4495, 15) & to_signed(1098457, 22)),
    std_logic_vector(to_signed(-4486, 15) & to_signed(1097335, 22)),
    std_logic_vector(to_signed(-4477, 15) & to_signed(1096214, 22)),
    std_logic_vector(to_signed(-4468, 15) & to_signed(1095096, 22)),
    std_logic_vector(to_signed(-4458, 15) & to_signed(1093980, 22)),
    std_logic_vector(to_signed(-4449, 15) & to_signed(1092867, 22)),
    std_logic_vector(to_signed(-4440, 15) & to_signed(1091756, 22)),
    std_logic_vector(to_signed(-4431, 15) & to_signed(1090647, 22)),
    std_logic_vector(to_signed(-4422, 15) & to_signed(1089540, 22)),
    std_logic_vector(to_signed(-4413, 15) & to_signed(1088436, 22)),
    std_logic_vector(to_signed(-4404, 15) & to_signed(1087333, 22)),
    std_logic_vector(to_signed(-4395, 15) & to_signed(1086234, 22)),
    std_logic_vector(to_signed(-4387, 15) & to_signed(1085136, 22)),
    std_logic_vector(to_signed(-4378, 15) & to_signed(1084040, 22)),
    std_logic_vector(to_signed(-4369, 15) & to_signed(1082947, 22)),
    std_logic_vector(to_signed(-4360, 15) & to_signed(1081856, 22)),
    std_logic_vector(to_signed(-4351, 15) & to_signed(1080767, 22)),
    std_logic_vector(to_signed(-4343, 15) & to_signed(1079680, 22)),
    std_logic_vector(to_signed(-4334, 15) & to_signed(1078596, 22)),
    std_logic_vector(to_signed(-4325, 15) & to_signed(1077513, 22)),
    std_logic_vector(to_signed(-4317, 15) & to_signed(1076433, 22)),
    std_logic_vector(to_signed(-4308, 15) & to_signed(1075355, 22)),
    std_logic_vector(to_signed(-4299, 15) & to_signed(1074279, 22)),
    std_logic_vector(to_signed(-4291, 15) & to_signed(1073205, 22)),
    std_logic_vector(to_signed(-4282, 15) & to_signed(1072134, 22)),
    std_logic_vector(to_signed(-4274, 15) & to_signed(1071064, 22)),
    std_logic_vector(to_signed(-4265, 15) & to_signed(1069997, 22)),
    std_logic_vector(to_signed(-4257, 15) & to_signed(1068932, 22)),
    std_logic_vector(to_signed(-4248, 15) & to_signed(1067869, 22)),
    std_logic_vector(to_signed(-4240, 15) & to_signed(1066808, 22)),
    std_logic_vector(to_signed(-4231, 15) & to_signed(1065749, 22)),
    std_logic_vector(to_signed(-4223, 15) & to_signed(1064692, 22)),
    std_logic_vector(to_signed(-4215, 15) & to_signed(1063637, 22)),
    std_logic_vector(to_signed(-4206, 15) & to_signed(1062585, 22)),
    std_logic_vector(to_signed(-4198, 15) & to_signed(1061534, 22)),
    std_logic_vector(to_signed(-4190, 15) & to_signed(1060486, 22)),
    std_logic_vector(to_signed(-4181, 15) & to_signed(1059439, 22)),
    std_logic_vector(to_signed(-4173, 15) & to_signed(1058395, 22)),
    std_logic_vector(to_signed(-4165, 15) & to_signed(1057353, 22)),
    std_logic_vector(to_signed(-4157, 15) & to_signed(1056313, 22)),
    std_logic_vector(to_signed(-4148, 15) & to_signed(1055275, 22)),
    std_logic_vector(to_signed(-4140, 15) & to_signed(1054238, 22)),
    std_logic_vector(to_signed(-4132, 15) & to_signed(1053204, 22)),
    std_logic_vector(to_signed(-4124, 15) & to_signed(1052172, 22)),
    std_logic_vector(to_signed(-4116, 15) & to_signed(1051142, 22)),
    std_logic_vector(to_signed(-4108, 15) & to_signed(1050114, 22)),
    std_logic_vector(to_signed(-4100, 15) & to_signed(1049088, 22))
  );

  -- Signals
  signal TableAddr : std_logic_vector(log2ceil(TableSize_c) - 1 downto 0);
  signal TableData : std_logic_vector(TableWidth_c - 1 downto 0);

begin

  -- *** Calculation Unit ***
  i_calc : entity work.psi_fix_lin_approx_calc
    generic map(
      InFmt_g     => InFmt_c,
      OutFmt_g    => OutFmt_c,
      OffsFmt_g   => OffsFmt_c,
      GradFmt_g   => GradFmt_c,
      TableSize_g => TableSize_c
    )
    port map(
      -- Control Signals
      clk_i        => clk_i,
      rst_i        => rst_i,
      -- Input
      vld_i        => vld_i,
      dat_i        => dat_i,
      -- Output
      vld_o        => vld_o,
      dat_o        => dat_o,
      -- Table Interface
      addr_table_o => TableAddr,
      data_table_i => TableData
    );

  -- *** Table ***
  p_table : process(clk_i)
  begin
    if rising_edge(clk_i) then
      TableData <= Table_c(to_integer(unsigned(TableAddr)));
    end if;
  end process;

end rtl;
