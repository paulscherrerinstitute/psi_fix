------------------------------------------------------------------------------
-- Libraries
------------------------------------------------------------------------------
library ieee;
	use ieee.std_logic_1164.all;
	use ieee.numeric_std.all;
	
library psi_common;
	use work.psi_fix_pkg.all;
	use psi_common.psi_common_math_pkg.all;
	
------------------------------------------------------------------------------
-- Entity Declaration
------------------------------------------------------------------------------
entity psi_fix_lin_approx_sin18b_dual is
	port (
		-- Control Signals
		Clk			: in 	std_logic;
		Rst			: in 	std_logic;
		-- Input
		InVldA		: in	std_logic;
		InDataA		: in	std_logic_vector(20-1 downto 0);		-- Format (0, 0, 20)
		InVldB		: in	std_logic;
		InDataB		: in	std_logic_vector(20-1 downto 0);		-- Format (0, 0, 20)
		-- Output
		OutVldA		: out	std_logic;
		OutDataA	: out	std_logic_vector(18-1 downto 0);		-- Format (1, 0, 17)
		OutVldB		: out	std_logic;
		OutDataB	: out	std_logic_vector(18-1 downto 0)		-- Format (1, 0, 17)		
	);
end entity;

------------------------------------------------------------------------------
-- Architecture Declaration
------------------------------------------------------------------------------
architecture rtl of psi_fix_lin_approx_sin18b_dual is

	-- Constants
	constant InFmt_c		: PsiFixFmt_t		:= (0, 0, 20);
	constant OutFmt_c		: PsiFixFmt_t		:= (1, 0, 17);
	constant OffsFmt_c		: PsiFixFmt_t		:= (1, 0, 19);
	constant GradFmt_c		: PsiFixFmt_t		:= (1, 3, 8);
	constant TableSize_c	: integer			:= 2048;
	constant TableWidth_c	: integer			:= 32;
	
	-- Table	
	type Table_t is array(0 to TableSize_c-1) of std_logic_vector(TableWidth_c-1 downto 0);
	constant Table_c : Table_t := (
		std_logic_vector(to_signed(1608, 12) & to_signed(804, 20)),
		std_logic_vector(to_signed(1608, 12) & to_signed(2413, 20)),
		std_logic_vector(to_signed(1608, 12) & to_signed(4021, 20)),
		std_logic_vector(to_signed(1608, 12) & to_signed(5630, 20)),
		std_logic_vector(to_signed(1608, 12) & to_signed(7238, 20)),
		std_logic_vector(to_signed(1608, 12) & to_signed(8846, 20)),
		std_logic_vector(to_signed(1608, 12) & to_signed(10454, 20)),
		std_logic_vector(to_signed(1608, 12) & to_signed(12063, 20)),
		std_logic_vector(to_signed(1608, 12) & to_signed(13671, 20)),
		std_logic_vector(to_signed(1608, 12) & to_signed(15278, 20)),
		std_logic_vector(to_signed(1608, 12) & to_signed(16886, 20)),
		std_logic_vector(to_signed(1607, 12) & to_signed(18494, 20)),
		std_logic_vector(to_signed(1607, 12) & to_signed(20101, 20)),
		std_logic_vector(to_signed(1607, 12) & to_signed(21708, 20)),
		std_logic_vector(to_signed(1607, 12) & to_signed(23315, 20)),
		std_logic_vector(to_signed(1607, 12) & to_signed(24922, 20)),
		std_logic_vector(to_signed(1606, 12) & to_signed(26529, 20)),
		std_logic_vector(to_signed(1606, 12) & to_signed(28135, 20)),
		std_logic_vector(to_signed(1606, 12) & to_signed(29741, 20)),
		std_logic_vector(to_signed(1606, 12) & to_signed(31347, 20)),
		std_logic_vector(to_signed(1605, 12) & to_signed(32952, 20)),
		std_logic_vector(to_signed(1605, 12) & to_signed(34557, 20)),
		std_logic_vector(to_signed(1605, 12) & to_signed(36162, 20)),
		std_logic_vector(to_signed(1604, 12) & to_signed(37767, 20)),
		std_logic_vector(to_signed(1604, 12) & to_signed(39371, 20)),
		std_logic_vector(to_signed(1604, 12) & to_signed(40974, 20)),
		std_logic_vector(to_signed(1603, 12) & to_signed(42578, 20)),
		std_logic_vector(to_signed(1603, 12) & to_signed(44181, 20)),
		std_logic_vector(to_signed(1602, 12) & to_signed(45783, 20)),
		std_logic_vector(to_signed(1602, 12) & to_signed(47386, 20)),
		std_logic_vector(to_signed(1601, 12) & to_signed(48987, 20)),
		std_logic_vector(to_signed(1601, 12) & to_signed(50588, 20)),
		std_logic_vector(to_signed(1600, 12) & to_signed(52189, 20)),
		std_logic_vector(to_signed(1600, 12) & to_signed(53789, 20)),
		std_logic_vector(to_signed(1599, 12) & to_signed(55389, 20)),
		std_logic_vector(to_signed(1599, 12) & to_signed(56988, 20)),
		std_logic_vector(to_signed(1598, 12) & to_signed(58587, 20)),
		std_logic_vector(to_signed(1598, 12) & to_signed(60185, 20)),
		std_logic_vector(to_signed(1597, 12) & to_signed(61783, 20)),
		std_logic_vector(to_signed(1597, 12) & to_signed(63380, 20)),
		std_logic_vector(to_signed(1596, 12) & to_signed(64976, 20)),
		std_logic_vector(to_signed(1595, 12) & to_signed(66572, 20)),
		std_logic_vector(to_signed(1595, 12) & to_signed(68167, 20)),
		std_logic_vector(to_signed(1594, 12) & to_signed(69762, 20)),
		std_logic_vector(to_signed(1594, 12) & to_signed(71355, 20)),
		std_logic_vector(to_signed(1593, 12) & to_signed(72949, 20)),
		std_logic_vector(to_signed(1592, 12) & to_signed(74541, 20)),
		std_logic_vector(to_signed(1591, 12) & to_signed(76133, 20)),
		std_logic_vector(to_signed(1591, 12) & to_signed(77724, 20)),
		std_logic_vector(to_signed(1590, 12) & to_signed(79314, 20)),
		std_logic_vector(to_signed(1589, 12) & to_signed(80904, 20)),
		std_logic_vector(to_signed(1588, 12) & to_signed(82493, 20)),
		std_logic_vector(to_signed(1588, 12) & to_signed(84081, 20)),
		std_logic_vector(to_signed(1587, 12) & to_signed(85668, 20)),
		std_logic_vector(to_signed(1586, 12) & to_signed(87254, 20)),
		std_logic_vector(to_signed(1585, 12) & to_signed(88840, 20)),
		std_logic_vector(to_signed(1584, 12) & to_signed(90425, 20)),
		std_logic_vector(to_signed(1584, 12) & to_signed(92009, 20)),
		std_logic_vector(to_signed(1583, 12) & to_signed(93592, 20)),
		std_logic_vector(to_signed(1582, 12) & to_signed(95174, 20)),
		std_logic_vector(to_signed(1581, 12) & to_signed(96755, 20)),
		std_logic_vector(to_signed(1580, 12) & to_signed(98336, 20)),
		std_logic_vector(to_signed(1579, 12) & to_signed(99915, 20)),
		std_logic_vector(to_signed(1578, 12) & to_signed(101494, 20)),
		std_logic_vector(to_signed(1577, 12) & to_signed(103071, 20)),
		std_logic_vector(to_signed(1576, 12) & to_signed(104648, 20)),
		std_logic_vector(to_signed(1575, 12) & to_signed(106224, 20)),
		std_logic_vector(to_signed(1574, 12) & to_signed(107798, 20)),
		std_logic_vector(to_signed(1573, 12) & to_signed(109372, 20)),
		std_logic_vector(to_signed(1572, 12) & to_signed(110944, 20)),
		std_logic_vector(to_signed(1571, 12) & to_signed(112516, 20)),
		std_logic_vector(to_signed(1570, 12) & to_signed(114086, 20)),
		std_logic_vector(to_signed(1569, 12) & to_signed(115656, 20)),
		std_logic_vector(to_signed(1568, 12) & to_signed(117224, 20)),
		std_logic_vector(to_signed(1567, 12) & to_signed(118791, 20)),
		std_logic_vector(to_signed(1566, 12) & to_signed(120357, 20)),
		std_logic_vector(to_signed(1564, 12) & to_signed(121922, 20)),
		std_logic_vector(to_signed(1563, 12) & to_signed(123486, 20)),
		std_logic_vector(to_signed(1562, 12) & to_signed(125049, 20)),
		std_logic_vector(to_signed(1561, 12) & to_signed(126610, 20)),
		std_logic_vector(to_signed(1560, 12) & to_signed(128171, 20)),
		std_logic_vector(to_signed(1558, 12) & to_signed(129730, 20)),
		std_logic_vector(to_signed(1557, 12) & to_signed(131288, 20)),
		std_logic_vector(to_signed(1556, 12) & to_signed(132844, 20)),
		std_logic_vector(to_signed(1555, 12) & to_signed(134400, 20)),
		std_logic_vector(to_signed(1553, 12) & to_signed(135954, 20)),
		std_logic_vector(to_signed(1552, 12) & to_signed(137506, 20)),
		std_logic_vector(to_signed(1551, 12) & to_signed(139058, 20)),
		std_logic_vector(to_signed(1550, 12) & to_signed(140608, 20)),
		std_logic_vector(to_signed(1548, 12) & to_signed(142157, 20)),
		std_logic_vector(to_signed(1547, 12) & to_signed(143705, 20)),
		std_logic_vector(to_signed(1546, 12) & to_signed(145251, 20)),
		std_logic_vector(to_signed(1544, 12) & to_signed(146796, 20)),
		std_logic_vector(to_signed(1543, 12) & to_signed(148339, 20)),
		std_logic_vector(to_signed(1541, 12) & to_signed(149881, 20)),
		std_logic_vector(to_signed(1540, 12) & to_signed(151422, 20)),
		std_logic_vector(to_signed(1539, 12) & to_signed(152961, 20)),
		std_logic_vector(to_signed(1537, 12) & to_signed(154499, 20)),
		std_logic_vector(to_signed(1536, 12) & to_signed(156035, 20)),
		std_logic_vector(to_signed(1534, 12) & to_signed(157570, 20)),
		std_logic_vector(to_signed(1533, 12) & to_signed(159103, 20)),
		std_logic_vector(to_signed(1531, 12) & to_signed(160635, 20)),
		std_logic_vector(to_signed(1530, 12) & to_signed(162166, 20)),
		std_logic_vector(to_signed(1528, 12) & to_signed(163694, 20)),
		std_logic_vector(to_signed(1527, 12) & to_signed(165222, 20)),
		std_logic_vector(to_signed(1525, 12) & to_signed(166748, 20)),
		std_logic_vector(to_signed(1523, 12) & to_signed(168272, 20)),
		std_logic_vector(to_signed(1522, 12) & to_signed(169794, 20)),
		std_logic_vector(to_signed(1520, 12) & to_signed(171315, 20)),
		std_logic_vector(to_signed(1519, 12) & to_signed(172835, 20)),
		std_logic_vector(to_signed(1517, 12) & to_signed(174352, 20)),
		std_logic_vector(to_signed(1515, 12) & to_signed(175869, 20)),
		std_logic_vector(to_signed(1514, 12) & to_signed(177383, 20)),
		std_logic_vector(to_signed(1512, 12) & to_signed(178896, 20)),
		std_logic_vector(to_signed(1510, 12) & to_signed(180407, 20)),
		std_logic_vector(to_signed(1509, 12) & to_signed(181916, 20)),
		std_logic_vector(to_signed(1507, 12) & to_signed(183424, 20)),
		std_logic_vector(to_signed(1505, 12) & to_signed(184930, 20)),
		std_logic_vector(to_signed(1503, 12) & to_signed(186434, 20)),
		std_logic_vector(to_signed(1502, 12) & to_signed(187937, 20)),
		std_logic_vector(to_signed(1500, 12) & to_signed(189437, 20)),
		std_logic_vector(to_signed(1498, 12) & to_signed(190936, 20)),
		std_logic_vector(to_signed(1496, 12) & to_signed(192433, 20)),
		std_logic_vector(to_signed(1494, 12) & to_signed(193929, 20)),
		std_logic_vector(to_signed(1493, 12) & to_signed(195422, 20)),
		std_logic_vector(to_signed(1491, 12) & to_signed(196914, 20)),
		std_logic_vector(to_signed(1489, 12) & to_signed(198404, 20)),
		std_logic_vector(to_signed(1487, 12) & to_signed(199892, 20)),
		std_logic_vector(to_signed(1485, 12) & to_signed(201378, 20)),
		std_logic_vector(to_signed(1483, 12) & to_signed(202862, 20)),
		std_logic_vector(to_signed(1481, 12) & to_signed(204344, 20)),
		std_logic_vector(to_signed(1479, 12) & to_signed(205824, 20)),
		std_logic_vector(to_signed(1477, 12) & to_signed(207303, 20)),
		std_logic_vector(to_signed(1475, 12) & to_signed(208779, 20)),
		std_logic_vector(to_signed(1473, 12) & to_signed(210254, 20)),
		std_logic_vector(to_signed(1471, 12) & to_signed(211726, 20)),
		std_logic_vector(to_signed(1469, 12) & to_signed(213197, 20)),
		std_logic_vector(to_signed(1467, 12) & to_signed(214665, 20)),
		std_logic_vector(to_signed(1465, 12) & to_signed(216131, 20)),
		std_logic_vector(to_signed(1463, 12) & to_signed(217596, 20)),
		std_logic_vector(to_signed(1461, 12) & to_signed(219058, 20)),
		std_logic_vector(to_signed(1459, 12) & to_signed(220519, 20)),
		std_logic_vector(to_signed(1457, 12) & to_signed(221977, 20)),
		std_logic_vector(to_signed(1455, 12) & to_signed(223433, 20)),
		std_logic_vector(to_signed(1453, 12) & to_signed(224887, 20)),
		std_logic_vector(to_signed(1451, 12) & to_signed(226339, 20)),
		std_logic_vector(to_signed(1449, 12) & to_signed(227789, 20)),
		std_logic_vector(to_signed(1447, 12) & to_signed(229236, 20)),
		std_logic_vector(to_signed(1444, 12) & to_signed(230682, 20)),
		std_logic_vector(to_signed(1442, 12) & to_signed(232125, 20)),
		std_logic_vector(to_signed(1440, 12) & to_signed(233566, 20)),
		std_logic_vector(to_signed(1438, 12) & to_signed(235005, 20)),
		std_logic_vector(to_signed(1436, 12) & to_signed(236442, 20)),
		std_logic_vector(to_signed(1433, 12) & to_signed(237877, 20)),
		std_logic_vector(to_signed(1431, 12) & to_signed(239309, 20)),
		std_logic_vector(to_signed(1429, 12) & to_signed(240739, 20)),
		std_logic_vector(to_signed(1427, 12) & to_signed(242167, 20)),
		std_logic_vector(to_signed(1424, 12) & to_signed(243592, 20)),
		std_logic_vector(to_signed(1422, 12) & to_signed(245015, 20)),
		std_logic_vector(to_signed(1420, 12) & to_signed(246436, 20)),
		std_logic_vector(to_signed(1417, 12) & to_signed(247855, 20)),
		std_logic_vector(to_signed(1415, 12) & to_signed(249271, 20)),
		std_logic_vector(to_signed(1413, 12) & to_signed(250685, 20)),
		std_logic_vector(to_signed(1410, 12) & to_signed(252096, 20)),
		std_logic_vector(to_signed(1408, 12) & to_signed(253506, 20)),
		std_logic_vector(to_signed(1406, 12) & to_signed(254912, 20)),
		std_logic_vector(to_signed(1403, 12) & to_signed(256317, 20)),
		std_logic_vector(to_signed(1401, 12) & to_signed(257719, 20)),
		std_logic_vector(to_signed(1398, 12) & to_signed(259118, 20)),
		std_logic_vector(to_signed(1396, 12) & to_signed(260515, 20)),
		std_logic_vector(to_signed(1393, 12) & to_signed(261910, 20)),
		std_logic_vector(to_signed(1391, 12) & to_signed(263302, 20)),
		std_logic_vector(to_signed(1388, 12) & to_signed(264692, 20)),
		std_logic_vector(to_signed(1386, 12) & to_signed(266079, 20)),
		std_logic_vector(to_signed(1383, 12) & to_signed(267464, 20)),
		std_logic_vector(to_signed(1381, 12) & to_signed(268846, 20)),
		std_logic_vector(to_signed(1378, 12) & to_signed(270225, 20)),
		std_logic_vector(to_signed(1376, 12) & to_signed(271602, 20)),
		std_logic_vector(to_signed(1373, 12) & to_signed(272977, 20)),
		std_logic_vector(to_signed(1371, 12) & to_signed(274349, 20)),
		std_logic_vector(to_signed(1368, 12) & to_signed(275718, 20)),
		std_logic_vector(to_signed(1365, 12) & to_signed(277085, 20)),
		std_logic_vector(to_signed(1363, 12) & to_signed(278449, 20)),
		std_logic_vector(to_signed(1360, 12) & to_signed(279811, 20)),
		std_logic_vector(to_signed(1358, 12) & to_signed(281170, 20)),
		std_logic_vector(to_signed(1355, 12) & to_signed(282526, 20)),
		std_logic_vector(to_signed(1352, 12) & to_signed(283880, 20)),
		std_logic_vector(to_signed(1350, 12) & to_signed(285231, 20)),
		std_logic_vector(to_signed(1347, 12) & to_signed(286579, 20)),
		std_logic_vector(to_signed(1344, 12) & to_signed(287925, 20)),
		std_logic_vector(to_signed(1342, 12) & to_signed(289267, 20)),
		std_logic_vector(to_signed(1339, 12) & to_signed(290608, 20)),
		std_logic_vector(to_signed(1336, 12) & to_signed(291945, 20)),
		std_logic_vector(to_signed(1333, 12) & to_signed(293280, 20)),
		std_logic_vector(to_signed(1331, 12) & to_signed(294611, 20)),
		std_logic_vector(to_signed(1328, 12) & to_signed(295941, 20)),
		std_logic_vector(to_signed(1325, 12) & to_signed(297267, 20)),
		std_logic_vector(to_signed(1322, 12) & to_signed(298590, 20)),
		std_logic_vector(to_signed(1319, 12) & to_signed(299911, 20)),
		std_logic_vector(to_signed(1316, 12) & to_signed(301229, 20)),
		std_logic_vector(to_signed(1314, 12) & to_signed(302544, 20)),
		std_logic_vector(to_signed(1311, 12) & to_signed(303856, 20)),
		std_logic_vector(to_signed(1308, 12) & to_signed(305166, 20)),
		std_logic_vector(to_signed(1305, 12) & to_signed(306472, 20)),
		std_logic_vector(to_signed(1302, 12) & to_signed(307776, 20)),
		std_logic_vector(to_signed(1299, 12) & to_signed(309077, 20)),
		std_logic_vector(to_signed(1296, 12) & to_signed(310374, 20)),
		std_logic_vector(to_signed(1293, 12) & to_signed(311669, 20)),
		std_logic_vector(to_signed(1290, 12) & to_signed(312961, 20)),
		std_logic_vector(to_signed(1288, 12) & to_signed(314250, 20)),
		std_logic_vector(to_signed(1285, 12) & to_signed(315536, 20)),
		std_logic_vector(to_signed(1282, 12) & to_signed(316819, 20)),
		std_logic_vector(to_signed(1279, 12) & to_signed(318099, 20)),
		std_logic_vector(to_signed(1276, 12) & to_signed(319377, 20)),
		std_logic_vector(to_signed(1273, 12) & to_signed(320651, 20)),
		std_logic_vector(to_signed(1270, 12) & to_signed(321922, 20)),
		std_logic_vector(to_signed(1267, 12) & to_signed(323190, 20)),
		std_logic_vector(to_signed(1263, 12) & to_signed(324455, 20)),
		std_logic_vector(to_signed(1260, 12) & to_signed(325717, 20)),
		std_logic_vector(to_signed(1257, 12) & to_signed(326976, 20)),
		std_logic_vector(to_signed(1254, 12) & to_signed(328231, 20)),
		std_logic_vector(to_signed(1251, 12) & to_signed(329484, 20)),
		std_logic_vector(to_signed(1248, 12) & to_signed(330734, 20)),
		std_logic_vector(to_signed(1245, 12) & to_signed(331980, 20)),
		std_logic_vector(to_signed(1242, 12) & to_signed(333224, 20)),
		std_logic_vector(to_signed(1239, 12) & to_signed(334464, 20)),
		std_logic_vector(to_signed(1236, 12) & to_signed(335701, 20)),
		std_logic_vector(to_signed(1232, 12) & to_signed(336935, 20)),
		std_logic_vector(to_signed(1229, 12) & to_signed(338166, 20)),
		std_logic_vector(to_signed(1226, 12) & to_signed(339393, 20)),
		std_logic_vector(to_signed(1223, 12) & to_signed(340618, 20)),
		std_logic_vector(to_signed(1220, 12) & to_signed(341839, 20)),
		std_logic_vector(to_signed(1216, 12) & to_signed(343057, 20)),
		std_logic_vector(to_signed(1213, 12) & to_signed(344271, 20)),
		std_logic_vector(to_signed(1210, 12) & to_signed(345483, 20)),
		std_logic_vector(to_signed(1207, 12) & to_signed(346691, 20)),
		std_logic_vector(to_signed(1203, 12) & to_signed(347896, 20)),
		std_logic_vector(to_signed(1200, 12) & to_signed(349098, 20)),
		std_logic_vector(to_signed(1197, 12) & to_signed(350296, 20)),
		std_logic_vector(to_signed(1193, 12) & to_signed(351491, 20)),
		std_logic_vector(to_signed(1190, 12) & to_signed(352683, 20)),
		std_logic_vector(to_signed(1187, 12) & to_signed(353872, 20)),
		std_logic_vector(to_signed(1183, 12) & to_signed(355057, 20)),
		std_logic_vector(to_signed(1180, 12) & to_signed(356239, 20)),
		std_logic_vector(to_signed(1177, 12) & to_signed(357417, 20)),
		std_logic_vector(to_signed(1173, 12) & to_signed(358592, 20)),
		std_logic_vector(to_signed(1170, 12) & to_signed(359764, 20)),
		std_logic_vector(to_signed(1167, 12) & to_signed(360932, 20)),
		std_logic_vector(to_signed(1163, 12) & to_signed(362097, 20)),
		std_logic_vector(to_signed(1160, 12) & to_signed(363259, 20)),
		std_logic_vector(to_signed(1156, 12) & to_signed(364417, 20)),
		std_logic_vector(to_signed(1153, 12) & to_signed(365571, 20)),
		std_logic_vector(to_signed(1150, 12) & to_signed(366723, 20)),
		std_logic_vector(to_signed(1146, 12) & to_signed(367870, 20)),
		std_logic_vector(to_signed(1143, 12) & to_signed(369015, 20)),
		std_logic_vector(to_signed(1139, 12) & to_signed(370156, 20)),
		std_logic_vector(to_signed(1136, 12) & to_signed(371293, 20)),
		std_logic_vector(to_signed(1132, 12) & to_signed(372427, 20)),
		std_logic_vector(to_signed(1129, 12) & to_signed(373557, 20)),
		std_logic_vector(to_signed(1125, 12) & to_signed(374684, 20)),
		std_logic_vector(to_signed(1122, 12) & to_signed(375807, 20)),
		std_logic_vector(to_signed(1118, 12) & to_signed(376927, 20)),
		std_logic_vector(to_signed(1114, 12) & to_signed(378043, 20)),
		std_logic_vector(to_signed(1111, 12) & to_signed(379156, 20)),
		std_logic_vector(to_signed(1107, 12) & to_signed(380265, 20)),
		std_logic_vector(to_signed(1104, 12) & to_signed(381371, 20)),
		std_logic_vector(to_signed(1100, 12) & to_signed(382473, 20)),
		std_logic_vector(to_signed(1097, 12) & to_signed(383571, 20)),
		std_logic_vector(to_signed(1093, 12) & to_signed(384666, 20)),
		std_logic_vector(to_signed(1089, 12) & to_signed(385757, 20)),
		std_logic_vector(to_signed(1086, 12) & to_signed(386844, 20)),
		std_logic_vector(to_signed(1082, 12) & to_signed(387928, 20)),
		std_logic_vector(to_signed(1078, 12) & to_signed(389008, 20)),
		std_logic_vector(to_signed(1075, 12) & to_signed(390085, 20)),
		std_logic_vector(to_signed(1071, 12) & to_signed(391158, 20)),
		std_logic_vector(to_signed(1067, 12) & to_signed(392227, 20)),
		std_logic_vector(to_signed(1064, 12) & to_signed(393293, 20)),
		std_logic_vector(to_signed(1060, 12) & to_signed(394354, 20)),
		std_logic_vector(to_signed(1056, 12) & to_signed(395412, 20)),
		std_logic_vector(to_signed(1052, 12) & to_signed(396467, 20)),
		std_logic_vector(to_signed(1049, 12) & to_signed(397517, 20)),
		std_logic_vector(to_signed(1045, 12) & to_signed(398564, 20)),
		std_logic_vector(to_signed(1041, 12) & to_signed(399607, 20)),
		std_logic_vector(to_signed(1037, 12) & to_signed(400647, 20)),
		std_logic_vector(to_signed(1034, 12) & to_signed(401682, 20)),
		std_logic_vector(to_signed(1030, 12) & to_signed(402714, 20)),
		std_logic_vector(to_signed(1026, 12) & to_signed(403742, 20)),
		std_logic_vector(to_signed(1022, 12) & to_signed(404766, 20)),
		std_logic_vector(to_signed(1019, 12) & to_signed(405787, 20)),
		std_logic_vector(to_signed(1015, 12) & to_signed(406803, 20)),
		std_logic_vector(to_signed(1011, 12) & to_signed(407816, 20)),
		std_logic_vector(to_signed(1007, 12) & to_signed(408825, 20)),
		std_logic_vector(to_signed(1003, 12) & to_signed(409830, 20)),
		std_logic_vector(to_signed(999, 12) & to_signed(410831, 20)),
		std_logic_vector(to_signed(995, 12) & to_signed(411829, 20)),
		std_logic_vector(to_signed(992, 12) & to_signed(412822, 20)),
		std_logic_vector(to_signed(988, 12) & to_signed(413812, 20)),
		std_logic_vector(to_signed(984, 12) & to_signed(414797, 20)),
		std_logic_vector(to_signed(980, 12) & to_signed(415779, 20)),
		std_logic_vector(to_signed(976, 12) & to_signed(416757, 20)),
		std_logic_vector(to_signed(972, 12) & to_signed(417731, 20)),
		std_logic_vector(to_signed(968, 12) & to_signed(418701, 20)),
		std_logic_vector(to_signed(964, 12) & to_signed(419667, 20)),
		std_logic_vector(to_signed(960, 12) & to_signed(420629, 20)),
		std_logic_vector(to_signed(956, 12) & to_signed(421587, 20)),
		std_logic_vector(to_signed(952, 12) & to_signed(422542, 20)),
		std_logic_vector(to_signed(948, 12) & to_signed(423492, 20)),
		std_logic_vector(to_signed(944, 12) & to_signed(424438, 20)),
		std_logic_vector(to_signed(940, 12) & to_signed(425380, 20)),
		std_logic_vector(to_signed(936, 12) & to_signed(426319, 20)),
		std_logic_vector(to_signed(932, 12) & to_signed(427253, 20)),
		std_logic_vector(to_signed(928, 12) & to_signed(428183, 20)),
		std_logic_vector(to_signed(924, 12) & to_signed(429109, 20)),
		std_logic_vector(to_signed(920, 12) & to_signed(430031, 20)),
		std_logic_vector(to_signed(916, 12) & to_signed(430949, 20)),
		std_logic_vector(to_signed(912, 12) & to_signed(431863, 20)),
		std_logic_vector(to_signed(908, 12) & to_signed(432773, 20)),
		std_logic_vector(to_signed(904, 12) & to_signed(433679, 20)),
		std_logic_vector(to_signed(900, 12) & to_signed(434581, 20)),
		std_logic_vector(to_signed(896, 12) & to_signed(435479, 20)),
		std_logic_vector(to_signed(892, 12) & to_signed(436373, 20)),
		std_logic_vector(to_signed(887, 12) & to_signed(437262, 20)),
		std_logic_vector(to_signed(883, 12) & to_signed(438147, 20)),
		std_logic_vector(to_signed(879, 12) & to_signed(439029, 20)),
		std_logic_vector(to_signed(875, 12) & to_signed(439906, 20)),
		std_logic_vector(to_signed(871, 12) & to_signed(440779, 20)),
		std_logic_vector(to_signed(867, 12) & to_signed(441648, 20)),
		std_logic_vector(to_signed(863, 12) & to_signed(442512, 20)),
		std_logic_vector(to_signed(858, 12) & to_signed(443373, 20)),
		std_logic_vector(to_signed(854, 12) & to_signed(444229, 20)),
		std_logic_vector(to_signed(850, 12) & to_signed(445081, 20)),
		std_logic_vector(to_signed(846, 12) & to_signed(445929, 20)),
		std_logic_vector(to_signed(842, 12) & to_signed(446773, 20)),
		std_logic_vector(to_signed(837, 12) & to_signed(447613, 20)),
		std_logic_vector(to_signed(833, 12) & to_signed(448448, 20)),
		std_logic_vector(to_signed(829, 12) & to_signed(449279, 20)),
		std_logic_vector(to_signed(825, 12) & to_signed(450106, 20)),
		std_logic_vector(to_signed(821, 12) & to_signed(450929, 20)),
		std_logic_vector(to_signed(816, 12) & to_signed(451747, 20)),
		std_logic_vector(to_signed(812, 12) & to_signed(452562, 20)),
		std_logic_vector(to_signed(808, 12) & to_signed(453372, 20)),
		std_logic_vector(to_signed(804, 12) & to_signed(454177, 20)),
		std_logic_vector(to_signed(799, 12) & to_signed(454979, 20)),
		std_logic_vector(to_signed(795, 12) & to_signed(455776, 20)),
		std_logic_vector(to_signed(791, 12) & to_signed(456569, 20)),
		std_logic_vector(to_signed(786, 12) & to_signed(457357, 20)),
		std_logic_vector(to_signed(782, 12) & to_signed(458141, 20)),
		std_logic_vector(to_signed(778, 12) & to_signed(458921, 20)),
		std_logic_vector(to_signed(773, 12) & to_signed(459697, 20)),
		std_logic_vector(to_signed(769, 12) & to_signed(460468, 20)),
		std_logic_vector(to_signed(765, 12) & to_signed(461235, 20)),
		std_logic_vector(to_signed(760, 12) & to_signed(461998, 20)),
		std_logic_vector(to_signed(756, 12) & to_signed(462756, 20)),
		std_logic_vector(to_signed(752, 12) & to_signed(463510, 20)),
		std_logic_vector(to_signed(747, 12) & to_signed(464259, 20)),
		std_logic_vector(to_signed(743, 12) & to_signed(465004, 20)),
		std_logic_vector(to_signed(739, 12) & to_signed(465745, 20)),
		std_logic_vector(to_signed(734, 12) & to_signed(466481, 20)),
		std_logic_vector(to_signed(730, 12) & to_signed(467213, 20)),
		std_logic_vector(to_signed(725, 12) & to_signed(467941, 20)),
		std_logic_vector(to_signed(721, 12) & to_signed(468664, 20)),
		std_logic_vector(to_signed(717, 12) & to_signed(469383, 20)),
		std_logic_vector(to_signed(712, 12) & to_signed(470097, 20)),
		std_logic_vector(to_signed(708, 12) & to_signed(470807, 20)),
		std_logic_vector(to_signed(703, 12) & to_signed(471513, 20)),
		std_logic_vector(to_signed(699, 12) & to_signed(472214, 20)),
		std_logic_vector(to_signed(694, 12) & to_signed(472911, 20)),
		std_logic_vector(to_signed(690, 12) & to_signed(473603, 20)),
		std_logic_vector(to_signed(685, 12) & to_signed(474290, 20)),
		std_logic_vector(to_signed(681, 12) & to_signed(474974, 20)),
		std_logic_vector(to_signed(677, 12) & to_signed(475652, 20)),
		std_logic_vector(to_signed(672, 12) & to_signed(476327, 20)),
		std_logic_vector(to_signed(668, 12) & to_signed(476997, 20)),
		std_logic_vector(to_signed(663, 12) & to_signed(477662, 20)),
		std_logic_vector(to_signed(659, 12) & to_signed(478323, 20)),
		std_logic_vector(to_signed(654, 12) & to_signed(478979, 20)),
		std_logic_vector(to_signed(650, 12) & to_signed(479631, 20)),
		std_logic_vector(to_signed(645, 12) & to_signed(480278, 20)),
		std_logic_vector(to_signed(641, 12) & to_signed(480921, 20)),
		std_logic_vector(to_signed(636, 12) & to_signed(481559, 20)),
		std_logic_vector(to_signed(631, 12) & to_signed(482193, 20)),
		std_logic_vector(to_signed(627, 12) & to_signed(482822, 20)),
		std_logic_vector(to_signed(622, 12) & to_signed(483447, 20)),
		std_logic_vector(to_signed(618, 12) & to_signed(484067, 20)),
		std_logic_vector(to_signed(613, 12) & to_signed(484682, 20)),
		std_logic_vector(to_signed(609, 12) & to_signed(485293, 20)),
		std_logic_vector(to_signed(604, 12) & to_signed(485900, 20)),
		std_logic_vector(to_signed(600, 12) & to_signed(486502, 20)),
		std_logic_vector(to_signed(595, 12) & to_signed(487099, 20)),
		std_logic_vector(to_signed(590, 12) & to_signed(487692, 20)),
		std_logic_vector(to_signed(586, 12) & to_signed(488280, 20)),
		std_logic_vector(to_signed(581, 12) & to_signed(488863, 20)),
		std_logic_vector(to_signed(577, 12) & to_signed(489442, 20)),
		std_logic_vector(to_signed(572, 12) & to_signed(490016, 20)),
		std_logic_vector(to_signed(567, 12) & to_signed(490586, 20)),
		std_logic_vector(to_signed(563, 12) & to_signed(491151, 20)),
		std_logic_vector(to_signed(558, 12) & to_signed(491711, 20)),
		std_logic_vector(to_signed(553, 12) & to_signed(492267, 20)),
		std_logic_vector(to_signed(549, 12) & to_signed(492818, 20)),
		std_logic_vector(to_signed(544, 12) & to_signed(493365, 20)),
		std_logic_vector(to_signed(540, 12) & to_signed(493907, 20)),
		std_logic_vector(to_signed(535, 12) & to_signed(494444, 20)),
		std_logic_vector(to_signed(530, 12) & to_signed(494977, 20)),
		std_logic_vector(to_signed(526, 12) & to_signed(495505, 20)),
		std_logic_vector(to_signed(521, 12) & to_signed(496028, 20)),
		std_logic_vector(to_signed(516, 12) & to_signed(496546, 20)),
		std_logic_vector(to_signed(512, 12) & to_signed(497060, 20)),
		std_logic_vector(to_signed(507, 12) & to_signed(497570, 20)),
		std_logic_vector(to_signed(502, 12) & to_signed(498074, 20)),
		std_logic_vector(to_signed(498, 12) & to_signed(498574, 20)),
		std_logic_vector(to_signed(493, 12) & to_signed(499069, 20)),
		std_logic_vector(to_signed(488, 12) & to_signed(499560, 20)),
		std_logic_vector(to_signed(483, 12) & to_signed(500045, 20)),
		std_logic_vector(to_signed(479, 12) & to_signed(500526, 20)),
		std_logic_vector(to_signed(474, 12) & to_signed(501003, 20)),
		std_logic_vector(to_signed(469, 12) & to_signed(501474, 20)),
		std_logic_vector(to_signed(465, 12) & to_signed(501941, 20)),
		std_logic_vector(to_signed(460, 12) & to_signed(502404, 20)),
		std_logic_vector(to_signed(455, 12) & to_signed(502861, 20)),
		std_logic_vector(to_signed(450, 12) & to_signed(503314, 20)),
		std_logic_vector(to_signed(446, 12) & to_signed(503762, 20)),
		std_logic_vector(to_signed(441, 12) & to_signed(504205, 20)),
		std_logic_vector(to_signed(436, 12) & to_signed(504644, 20)),
		std_logic_vector(to_signed(431, 12) & to_signed(505077, 20)),
		std_logic_vector(to_signed(427, 12) & to_signed(505506, 20)),
		std_logic_vector(to_signed(422, 12) & to_signed(505931, 20)),
		std_logic_vector(to_signed(417, 12) & to_signed(506350, 20)),
		std_logic_vector(to_signed(412, 12) & to_signed(506765, 20)),
		std_logic_vector(to_signed(408, 12) & to_signed(507175, 20)),
		std_logic_vector(to_signed(403, 12) & to_signed(507580, 20)),
		std_logic_vector(to_signed(398, 12) & to_signed(507980, 20)),
		std_logic_vector(to_signed(393, 12) & to_signed(508376, 20)),
		std_logic_vector(to_signed(388, 12) & to_signed(508767, 20)),
		std_logic_vector(to_signed(384, 12) & to_signed(509153, 20)),
		std_logic_vector(to_signed(379, 12) & to_signed(509534, 20)),
		std_logic_vector(to_signed(374, 12) & to_signed(509910, 20)),
		std_logic_vector(to_signed(369, 12) & to_signed(510282, 20)),
		std_logic_vector(to_signed(364, 12) & to_signed(510649, 20)),
		std_logic_vector(to_signed(360, 12) & to_signed(511011, 20)),
		std_logic_vector(to_signed(355, 12) & to_signed(511368, 20)),
		std_logic_vector(to_signed(350, 12) & to_signed(511721, 20)),
		std_logic_vector(to_signed(345, 12) & to_signed(512068, 20)),
		std_logic_vector(to_signed(340, 12) & to_signed(512411, 20)),
		std_logic_vector(to_signed(336, 12) & to_signed(512749, 20)),
		std_logic_vector(to_signed(331, 12) & to_signed(513082, 20)),
		std_logic_vector(to_signed(326, 12) & to_signed(513410, 20)),
		std_logic_vector(to_signed(321, 12) & to_signed(513734, 20)),
		std_logic_vector(to_signed(316, 12) & to_signed(514053, 20)),
		std_logic_vector(to_signed(311, 12) & to_signed(514366, 20)),
		std_logic_vector(to_signed(307, 12) & to_signed(514675, 20)),
		std_logic_vector(to_signed(302, 12) & to_signed(514979, 20)),
		std_logic_vector(to_signed(297, 12) & to_signed(515279, 20)),
		std_logic_vector(to_signed(292, 12) & to_signed(515573, 20)),
		std_logic_vector(to_signed(287, 12) & to_signed(515863, 20)),
		std_logic_vector(to_signed(282, 12) & to_signed(516147, 20)),
		std_logic_vector(to_signed(277, 12) & to_signed(516427, 20)),
		std_logic_vector(to_signed(273, 12) & to_signed(516702, 20)),
		std_logic_vector(to_signed(268, 12) & to_signed(516972, 20)),
		std_logic_vector(to_signed(263, 12) & to_signed(517238, 20)),
		std_logic_vector(to_signed(258, 12) & to_signed(517498, 20)),
		std_logic_vector(to_signed(253, 12) & to_signed(517753, 20)),
		std_logic_vector(to_signed(248, 12) & to_signed(518004, 20)),
		std_logic_vector(to_signed(243, 12) & to_signed(518250, 20)),
		std_logic_vector(to_signed(238, 12) & to_signed(518491, 20)),
		std_logic_vector(to_signed(234, 12) & to_signed(518727, 20)),
		std_logic_vector(to_signed(229, 12) & to_signed(518958, 20)),
		std_logic_vector(to_signed(224, 12) & to_signed(519184, 20)),
		std_logic_vector(to_signed(219, 12) & to_signed(519406, 20)),
		std_logic_vector(to_signed(214, 12) & to_signed(519622, 20)),
		std_logic_vector(to_signed(209, 12) & to_signed(519834, 20)),
		std_logic_vector(to_signed(204, 12) & to_signed(520040, 20)),
		std_logic_vector(to_signed(199, 12) & to_signed(520242, 20)),
		std_logic_vector(to_signed(194, 12) & to_signed(520439, 20)),
		std_logic_vector(to_signed(190, 12) & to_signed(520631, 20)),
		std_logic_vector(to_signed(185, 12) & to_signed(520818, 20)),
		std_logic_vector(to_signed(180, 12) & to_signed(521000, 20)),
		std_logic_vector(to_signed(175, 12) & to_signed(521178, 20)),
		std_logic_vector(to_signed(170, 12) & to_signed(521350, 20)),
		std_logic_vector(to_signed(165, 12) & to_signed(521517, 20)),
		std_logic_vector(to_signed(160, 12) & to_signed(521680, 20)),
		std_logic_vector(to_signed(155, 12) & to_signed(521838, 20)),
		std_logic_vector(to_signed(150, 12) & to_signed(521990, 20)),
		std_logic_vector(to_signed(145, 12) & to_signed(522138, 20)),
		std_logic_vector(to_signed(140, 12) & to_signed(522281, 20)),
		std_logic_vector(to_signed(136, 12) & to_signed(522419, 20)),
		std_logic_vector(to_signed(131, 12) & to_signed(522552, 20)),
		std_logic_vector(to_signed(126, 12) & to_signed(522680, 20)),
		std_logic_vector(to_signed(121, 12) & to_signed(522804, 20)),
		std_logic_vector(to_signed(116, 12) & to_signed(522922, 20)),
		std_logic_vector(to_signed(111, 12) & to_signed(523035, 20)),
		std_logic_vector(to_signed(106, 12) & to_signed(523144, 20)),
		std_logic_vector(to_signed(101, 12) & to_signed(523247, 20)),
		std_logic_vector(to_signed(96, 12) & to_signed(523346, 20)),
		std_logic_vector(to_signed(91, 12) & to_signed(523440, 20)),
		std_logic_vector(to_signed(86, 12) & to_signed(523529, 20)),
		std_logic_vector(to_signed(81, 12) & to_signed(523612, 20)),
		std_logic_vector(to_signed(76, 12) & to_signed(523691, 20)),
		std_logic_vector(to_signed(72, 12) & to_signed(523765, 20)),
		std_logic_vector(to_signed(67, 12) & to_signed(523834, 20)),
		std_logic_vector(to_signed(62, 12) & to_signed(523899, 20)),
		std_logic_vector(to_signed(57, 12) & to_signed(523958, 20)),
		std_logic_vector(to_signed(52, 12) & to_signed(524012, 20)),
		std_logic_vector(to_signed(47, 12) & to_signed(524061, 20)),
		std_logic_vector(to_signed(42, 12) & to_signed(524106, 20)),
		std_logic_vector(to_signed(37, 12) & to_signed(524145, 20)),
		std_logic_vector(to_signed(32, 12) & to_signed(524180, 20)),
		std_logic_vector(to_signed(27, 12) & to_signed(524209, 20)),
		std_logic_vector(to_signed(22, 12) & to_signed(524234, 20)),
		std_logic_vector(to_signed(17, 12) & to_signed(524254, 20)),
		std_logic_vector(to_signed(12, 12) & to_signed(524269, 20)),
		std_logic_vector(to_signed(7, 12) & to_signed(524278, 20)),
		std_logic_vector(to_signed(2, 12) & to_signed(524283, 20)),
		std_logic_vector(to_signed(-2, 12) & to_signed(524283, 20)),
		std_logic_vector(to_signed(-7, 12) & to_signed(524278, 20)),
		std_logic_vector(to_signed(-12, 12) & to_signed(524269, 20)),
		std_logic_vector(to_signed(-17, 12) & to_signed(524254, 20)),
		std_logic_vector(to_signed(-22, 12) & to_signed(524234, 20)),
		std_logic_vector(to_signed(-27, 12) & to_signed(524209, 20)),
		std_logic_vector(to_signed(-32, 12) & to_signed(524180, 20)),
		std_logic_vector(to_signed(-37, 12) & to_signed(524145, 20)),
		std_logic_vector(to_signed(-42, 12) & to_signed(524106, 20)),
		std_logic_vector(to_signed(-47, 12) & to_signed(524061, 20)),
		std_logic_vector(to_signed(-52, 12) & to_signed(524012, 20)),
		std_logic_vector(to_signed(-57, 12) & to_signed(523958, 20)),
		std_logic_vector(to_signed(-62, 12) & to_signed(523899, 20)),
		std_logic_vector(to_signed(-67, 12) & to_signed(523834, 20)),
		std_logic_vector(to_signed(-72, 12) & to_signed(523765, 20)),
		std_logic_vector(to_signed(-76, 12) & to_signed(523691, 20)),
		std_logic_vector(to_signed(-81, 12) & to_signed(523612, 20)),
		std_logic_vector(to_signed(-86, 12) & to_signed(523529, 20)),
		std_logic_vector(to_signed(-91, 12) & to_signed(523440, 20)),
		std_logic_vector(to_signed(-96, 12) & to_signed(523346, 20)),
		std_logic_vector(to_signed(-101, 12) & to_signed(523247, 20)),
		std_logic_vector(to_signed(-106, 12) & to_signed(523144, 20)),
		std_logic_vector(to_signed(-111, 12) & to_signed(523035, 20)),
		std_logic_vector(to_signed(-116, 12) & to_signed(522922, 20)),
		std_logic_vector(to_signed(-121, 12) & to_signed(522804, 20)),
		std_logic_vector(to_signed(-126, 12) & to_signed(522680, 20)),
		std_logic_vector(to_signed(-131, 12) & to_signed(522552, 20)),
		std_logic_vector(to_signed(-136, 12) & to_signed(522419, 20)),
		std_logic_vector(to_signed(-140, 12) & to_signed(522281, 20)),
		std_logic_vector(to_signed(-145, 12) & to_signed(522138, 20)),
		std_logic_vector(to_signed(-150, 12) & to_signed(521990, 20)),
		std_logic_vector(to_signed(-155, 12) & to_signed(521838, 20)),
		std_logic_vector(to_signed(-160, 12) & to_signed(521680, 20)),
		std_logic_vector(to_signed(-165, 12) & to_signed(521517, 20)),
		std_logic_vector(to_signed(-170, 12) & to_signed(521350, 20)),
		std_logic_vector(to_signed(-175, 12) & to_signed(521178, 20)),
		std_logic_vector(to_signed(-180, 12) & to_signed(521000, 20)),
		std_logic_vector(to_signed(-185, 12) & to_signed(520818, 20)),
		std_logic_vector(to_signed(-190, 12) & to_signed(520631, 20)),
		std_logic_vector(to_signed(-194, 12) & to_signed(520439, 20)),
		std_logic_vector(to_signed(-199, 12) & to_signed(520242, 20)),
		std_logic_vector(to_signed(-204, 12) & to_signed(520040, 20)),
		std_logic_vector(to_signed(-209, 12) & to_signed(519834, 20)),
		std_logic_vector(to_signed(-214, 12) & to_signed(519622, 20)),
		std_logic_vector(to_signed(-219, 12) & to_signed(519406, 20)),
		std_logic_vector(to_signed(-224, 12) & to_signed(519184, 20)),
		std_logic_vector(to_signed(-229, 12) & to_signed(518958, 20)),
		std_logic_vector(to_signed(-234, 12) & to_signed(518727, 20)),
		std_logic_vector(to_signed(-238, 12) & to_signed(518491, 20)),
		std_logic_vector(to_signed(-243, 12) & to_signed(518250, 20)),
		std_logic_vector(to_signed(-248, 12) & to_signed(518004, 20)),
		std_logic_vector(to_signed(-253, 12) & to_signed(517753, 20)),
		std_logic_vector(to_signed(-258, 12) & to_signed(517498, 20)),
		std_logic_vector(to_signed(-263, 12) & to_signed(517238, 20)),
		std_logic_vector(to_signed(-268, 12) & to_signed(516972, 20)),
		std_logic_vector(to_signed(-273, 12) & to_signed(516702, 20)),
		std_logic_vector(to_signed(-277, 12) & to_signed(516427, 20)),
		std_logic_vector(to_signed(-282, 12) & to_signed(516147, 20)),
		std_logic_vector(to_signed(-287, 12) & to_signed(515863, 20)),
		std_logic_vector(to_signed(-292, 12) & to_signed(515573, 20)),
		std_logic_vector(to_signed(-297, 12) & to_signed(515279, 20)),
		std_logic_vector(to_signed(-302, 12) & to_signed(514979, 20)),
		std_logic_vector(to_signed(-307, 12) & to_signed(514675, 20)),
		std_logic_vector(to_signed(-311, 12) & to_signed(514366, 20)),
		std_logic_vector(to_signed(-316, 12) & to_signed(514053, 20)),
		std_logic_vector(to_signed(-321, 12) & to_signed(513734, 20)),
		std_logic_vector(to_signed(-326, 12) & to_signed(513410, 20)),
		std_logic_vector(to_signed(-331, 12) & to_signed(513082, 20)),
		std_logic_vector(to_signed(-336, 12) & to_signed(512749, 20)),
		std_logic_vector(to_signed(-340, 12) & to_signed(512411, 20)),
		std_logic_vector(to_signed(-345, 12) & to_signed(512068, 20)),
		std_logic_vector(to_signed(-350, 12) & to_signed(511721, 20)),
		std_logic_vector(to_signed(-355, 12) & to_signed(511368, 20)),
		std_logic_vector(to_signed(-360, 12) & to_signed(511011, 20)),
		std_logic_vector(to_signed(-364, 12) & to_signed(510649, 20)),
		std_logic_vector(to_signed(-369, 12) & to_signed(510282, 20)),
		std_logic_vector(to_signed(-374, 12) & to_signed(509910, 20)),
		std_logic_vector(to_signed(-379, 12) & to_signed(509534, 20)),
		std_logic_vector(to_signed(-384, 12) & to_signed(509153, 20)),
		std_logic_vector(to_signed(-388, 12) & to_signed(508767, 20)),
		std_logic_vector(to_signed(-393, 12) & to_signed(508376, 20)),
		std_logic_vector(to_signed(-398, 12) & to_signed(507980, 20)),
		std_logic_vector(to_signed(-403, 12) & to_signed(507580, 20)),
		std_logic_vector(to_signed(-408, 12) & to_signed(507175, 20)),
		std_logic_vector(to_signed(-412, 12) & to_signed(506765, 20)),
		std_logic_vector(to_signed(-417, 12) & to_signed(506350, 20)),
		std_logic_vector(to_signed(-422, 12) & to_signed(505931, 20)),
		std_logic_vector(to_signed(-427, 12) & to_signed(505506, 20)),
		std_logic_vector(to_signed(-431, 12) & to_signed(505077, 20)),
		std_logic_vector(to_signed(-436, 12) & to_signed(504644, 20)),
		std_logic_vector(to_signed(-441, 12) & to_signed(504205, 20)),
		std_logic_vector(to_signed(-446, 12) & to_signed(503762, 20)),
		std_logic_vector(to_signed(-450, 12) & to_signed(503314, 20)),
		std_logic_vector(to_signed(-455, 12) & to_signed(502861, 20)),
		std_logic_vector(to_signed(-460, 12) & to_signed(502404, 20)),
		std_logic_vector(to_signed(-465, 12) & to_signed(501941, 20)),
		std_logic_vector(to_signed(-469, 12) & to_signed(501474, 20)),
		std_logic_vector(to_signed(-474, 12) & to_signed(501003, 20)),
		std_logic_vector(to_signed(-479, 12) & to_signed(500526, 20)),
		std_logic_vector(to_signed(-483, 12) & to_signed(500045, 20)),
		std_logic_vector(to_signed(-488, 12) & to_signed(499560, 20)),
		std_logic_vector(to_signed(-493, 12) & to_signed(499069, 20)),
		std_logic_vector(to_signed(-498, 12) & to_signed(498574, 20)),
		std_logic_vector(to_signed(-502, 12) & to_signed(498074, 20)),
		std_logic_vector(to_signed(-507, 12) & to_signed(497570, 20)),
		std_logic_vector(to_signed(-512, 12) & to_signed(497060, 20)),
		std_logic_vector(to_signed(-516, 12) & to_signed(496546, 20)),
		std_logic_vector(to_signed(-521, 12) & to_signed(496028, 20)),
		std_logic_vector(to_signed(-526, 12) & to_signed(495505, 20)),
		std_logic_vector(to_signed(-530, 12) & to_signed(494977, 20)),
		std_logic_vector(to_signed(-535, 12) & to_signed(494444, 20)),
		std_logic_vector(to_signed(-540, 12) & to_signed(493907, 20)),
		std_logic_vector(to_signed(-544, 12) & to_signed(493365, 20)),
		std_logic_vector(to_signed(-549, 12) & to_signed(492818, 20)),
		std_logic_vector(to_signed(-553, 12) & to_signed(492267, 20)),
		std_logic_vector(to_signed(-558, 12) & to_signed(491711, 20)),
		std_logic_vector(to_signed(-563, 12) & to_signed(491151, 20)),
		std_logic_vector(to_signed(-567, 12) & to_signed(490586, 20)),
		std_logic_vector(to_signed(-572, 12) & to_signed(490016, 20)),
		std_logic_vector(to_signed(-577, 12) & to_signed(489442, 20)),
		std_logic_vector(to_signed(-581, 12) & to_signed(488863, 20)),
		std_logic_vector(to_signed(-586, 12) & to_signed(488280, 20)),
		std_logic_vector(to_signed(-590, 12) & to_signed(487692, 20)),
		std_logic_vector(to_signed(-595, 12) & to_signed(487099, 20)),
		std_logic_vector(to_signed(-600, 12) & to_signed(486502, 20)),
		std_logic_vector(to_signed(-604, 12) & to_signed(485900, 20)),
		std_logic_vector(to_signed(-609, 12) & to_signed(485293, 20)),
		std_logic_vector(to_signed(-613, 12) & to_signed(484682, 20)),
		std_logic_vector(to_signed(-618, 12) & to_signed(484067, 20)),
		std_logic_vector(to_signed(-622, 12) & to_signed(483447, 20)),
		std_logic_vector(to_signed(-627, 12) & to_signed(482822, 20)),
		std_logic_vector(to_signed(-631, 12) & to_signed(482193, 20)),
		std_logic_vector(to_signed(-636, 12) & to_signed(481559, 20)),
		std_logic_vector(to_signed(-641, 12) & to_signed(480921, 20)),
		std_logic_vector(to_signed(-645, 12) & to_signed(480278, 20)),
		std_logic_vector(to_signed(-650, 12) & to_signed(479631, 20)),
		std_logic_vector(to_signed(-654, 12) & to_signed(478979, 20)),
		std_logic_vector(to_signed(-659, 12) & to_signed(478323, 20)),
		std_logic_vector(to_signed(-663, 12) & to_signed(477662, 20)),
		std_logic_vector(to_signed(-668, 12) & to_signed(476997, 20)),
		std_logic_vector(to_signed(-672, 12) & to_signed(476327, 20)),
		std_logic_vector(to_signed(-677, 12) & to_signed(475652, 20)),
		std_logic_vector(to_signed(-681, 12) & to_signed(474974, 20)),
		std_logic_vector(to_signed(-685, 12) & to_signed(474290, 20)),
		std_logic_vector(to_signed(-690, 12) & to_signed(473603, 20)),
		std_logic_vector(to_signed(-694, 12) & to_signed(472911, 20)),
		std_logic_vector(to_signed(-699, 12) & to_signed(472214, 20)),
		std_logic_vector(to_signed(-703, 12) & to_signed(471513, 20)),
		std_logic_vector(to_signed(-708, 12) & to_signed(470807, 20)),
		std_logic_vector(to_signed(-712, 12) & to_signed(470097, 20)),
		std_logic_vector(to_signed(-717, 12) & to_signed(469383, 20)),
		std_logic_vector(to_signed(-721, 12) & to_signed(468664, 20)),
		std_logic_vector(to_signed(-725, 12) & to_signed(467941, 20)),
		std_logic_vector(to_signed(-730, 12) & to_signed(467213, 20)),
		std_logic_vector(to_signed(-734, 12) & to_signed(466481, 20)),
		std_logic_vector(to_signed(-739, 12) & to_signed(465745, 20)),
		std_logic_vector(to_signed(-743, 12) & to_signed(465004, 20)),
		std_logic_vector(to_signed(-747, 12) & to_signed(464259, 20)),
		std_logic_vector(to_signed(-752, 12) & to_signed(463510, 20)),
		std_logic_vector(to_signed(-756, 12) & to_signed(462756, 20)),
		std_logic_vector(to_signed(-760, 12) & to_signed(461998, 20)),
		std_logic_vector(to_signed(-765, 12) & to_signed(461235, 20)),
		std_logic_vector(to_signed(-769, 12) & to_signed(460468, 20)),
		std_logic_vector(to_signed(-773, 12) & to_signed(459697, 20)),
		std_logic_vector(to_signed(-778, 12) & to_signed(458921, 20)),
		std_logic_vector(to_signed(-782, 12) & to_signed(458141, 20)),
		std_logic_vector(to_signed(-786, 12) & to_signed(457357, 20)),
		std_logic_vector(to_signed(-791, 12) & to_signed(456569, 20)),
		std_logic_vector(to_signed(-795, 12) & to_signed(455776, 20)),
		std_logic_vector(to_signed(-799, 12) & to_signed(454979, 20)),
		std_logic_vector(to_signed(-804, 12) & to_signed(454177, 20)),
		std_logic_vector(to_signed(-808, 12) & to_signed(453372, 20)),
		std_logic_vector(to_signed(-812, 12) & to_signed(452562, 20)),
		std_logic_vector(to_signed(-816, 12) & to_signed(451747, 20)),
		std_logic_vector(to_signed(-821, 12) & to_signed(450929, 20)),
		std_logic_vector(to_signed(-825, 12) & to_signed(450106, 20)),
		std_logic_vector(to_signed(-829, 12) & to_signed(449279, 20)),
		std_logic_vector(to_signed(-833, 12) & to_signed(448448, 20)),
		std_logic_vector(to_signed(-837, 12) & to_signed(447613, 20)),
		std_logic_vector(to_signed(-842, 12) & to_signed(446773, 20)),
		std_logic_vector(to_signed(-846, 12) & to_signed(445929, 20)),
		std_logic_vector(to_signed(-850, 12) & to_signed(445081, 20)),
		std_logic_vector(to_signed(-854, 12) & to_signed(444229, 20)),
		std_logic_vector(to_signed(-858, 12) & to_signed(443373, 20)),
		std_logic_vector(to_signed(-863, 12) & to_signed(442512, 20)),
		std_logic_vector(to_signed(-867, 12) & to_signed(441648, 20)),
		std_logic_vector(to_signed(-871, 12) & to_signed(440779, 20)),
		std_logic_vector(to_signed(-875, 12) & to_signed(439906, 20)),
		std_logic_vector(to_signed(-879, 12) & to_signed(439029, 20)),
		std_logic_vector(to_signed(-883, 12) & to_signed(438147, 20)),
		std_logic_vector(to_signed(-887, 12) & to_signed(437262, 20)),
		std_logic_vector(to_signed(-892, 12) & to_signed(436373, 20)),
		std_logic_vector(to_signed(-896, 12) & to_signed(435479, 20)),
		std_logic_vector(to_signed(-900, 12) & to_signed(434581, 20)),
		std_logic_vector(to_signed(-904, 12) & to_signed(433679, 20)),
		std_logic_vector(to_signed(-908, 12) & to_signed(432773, 20)),
		std_logic_vector(to_signed(-912, 12) & to_signed(431863, 20)),
		std_logic_vector(to_signed(-916, 12) & to_signed(430949, 20)),
		std_logic_vector(to_signed(-920, 12) & to_signed(430031, 20)),
		std_logic_vector(to_signed(-924, 12) & to_signed(429109, 20)),
		std_logic_vector(to_signed(-928, 12) & to_signed(428183, 20)),
		std_logic_vector(to_signed(-932, 12) & to_signed(427253, 20)),
		std_logic_vector(to_signed(-936, 12) & to_signed(426319, 20)),
		std_logic_vector(to_signed(-940, 12) & to_signed(425380, 20)),
		std_logic_vector(to_signed(-944, 12) & to_signed(424438, 20)),
		std_logic_vector(to_signed(-948, 12) & to_signed(423492, 20)),
		std_logic_vector(to_signed(-952, 12) & to_signed(422542, 20)),
		std_logic_vector(to_signed(-956, 12) & to_signed(421587, 20)),
		std_logic_vector(to_signed(-960, 12) & to_signed(420629, 20)),
		std_logic_vector(to_signed(-964, 12) & to_signed(419667, 20)),
		std_logic_vector(to_signed(-968, 12) & to_signed(418701, 20)),
		std_logic_vector(to_signed(-972, 12) & to_signed(417731, 20)),
		std_logic_vector(to_signed(-976, 12) & to_signed(416757, 20)),
		std_logic_vector(to_signed(-980, 12) & to_signed(415779, 20)),
		std_logic_vector(to_signed(-984, 12) & to_signed(414797, 20)),
		std_logic_vector(to_signed(-988, 12) & to_signed(413812, 20)),
		std_logic_vector(to_signed(-992, 12) & to_signed(412822, 20)),
		std_logic_vector(to_signed(-995, 12) & to_signed(411829, 20)),
		std_logic_vector(to_signed(-999, 12) & to_signed(410831, 20)),
		std_logic_vector(to_signed(-1003, 12) & to_signed(409830, 20)),
		std_logic_vector(to_signed(-1007, 12) & to_signed(408825, 20)),
		std_logic_vector(to_signed(-1011, 12) & to_signed(407816, 20)),
		std_logic_vector(to_signed(-1015, 12) & to_signed(406803, 20)),
		std_logic_vector(to_signed(-1019, 12) & to_signed(405787, 20)),
		std_logic_vector(to_signed(-1022, 12) & to_signed(404766, 20)),
		std_logic_vector(to_signed(-1026, 12) & to_signed(403742, 20)),
		std_logic_vector(to_signed(-1030, 12) & to_signed(402714, 20)),
		std_logic_vector(to_signed(-1034, 12) & to_signed(401682, 20)),
		std_logic_vector(to_signed(-1037, 12) & to_signed(400647, 20)),
		std_logic_vector(to_signed(-1041, 12) & to_signed(399607, 20)),
		std_logic_vector(to_signed(-1045, 12) & to_signed(398564, 20)),
		std_logic_vector(to_signed(-1049, 12) & to_signed(397517, 20)),
		std_logic_vector(to_signed(-1052, 12) & to_signed(396467, 20)),
		std_logic_vector(to_signed(-1056, 12) & to_signed(395412, 20)),
		std_logic_vector(to_signed(-1060, 12) & to_signed(394354, 20)),
		std_logic_vector(to_signed(-1064, 12) & to_signed(393293, 20)),
		std_logic_vector(to_signed(-1067, 12) & to_signed(392227, 20)),
		std_logic_vector(to_signed(-1071, 12) & to_signed(391158, 20)),
		std_logic_vector(to_signed(-1075, 12) & to_signed(390085, 20)),
		std_logic_vector(to_signed(-1078, 12) & to_signed(389008, 20)),
		std_logic_vector(to_signed(-1082, 12) & to_signed(387928, 20)),
		std_logic_vector(to_signed(-1086, 12) & to_signed(386844, 20)),
		std_logic_vector(to_signed(-1089, 12) & to_signed(385757, 20)),
		std_logic_vector(to_signed(-1093, 12) & to_signed(384666, 20)),
		std_logic_vector(to_signed(-1097, 12) & to_signed(383571, 20)),
		std_logic_vector(to_signed(-1100, 12) & to_signed(382473, 20)),
		std_logic_vector(to_signed(-1104, 12) & to_signed(381371, 20)),
		std_logic_vector(to_signed(-1107, 12) & to_signed(380265, 20)),
		std_logic_vector(to_signed(-1111, 12) & to_signed(379156, 20)),
		std_logic_vector(to_signed(-1114, 12) & to_signed(378043, 20)),
		std_logic_vector(to_signed(-1118, 12) & to_signed(376927, 20)),
		std_logic_vector(to_signed(-1122, 12) & to_signed(375807, 20)),
		std_logic_vector(to_signed(-1125, 12) & to_signed(374684, 20)),
		std_logic_vector(to_signed(-1129, 12) & to_signed(373557, 20)),
		std_logic_vector(to_signed(-1132, 12) & to_signed(372427, 20)),
		std_logic_vector(to_signed(-1136, 12) & to_signed(371293, 20)),
		std_logic_vector(to_signed(-1139, 12) & to_signed(370156, 20)),
		std_logic_vector(to_signed(-1143, 12) & to_signed(369015, 20)),
		std_logic_vector(to_signed(-1146, 12) & to_signed(367870, 20)),
		std_logic_vector(to_signed(-1150, 12) & to_signed(366723, 20)),
		std_logic_vector(to_signed(-1153, 12) & to_signed(365571, 20)),
		std_logic_vector(to_signed(-1156, 12) & to_signed(364417, 20)),
		std_logic_vector(to_signed(-1160, 12) & to_signed(363259, 20)),
		std_logic_vector(to_signed(-1163, 12) & to_signed(362097, 20)),
		std_logic_vector(to_signed(-1167, 12) & to_signed(360932, 20)),
		std_logic_vector(to_signed(-1170, 12) & to_signed(359764, 20)),
		std_logic_vector(to_signed(-1173, 12) & to_signed(358592, 20)),
		std_logic_vector(to_signed(-1177, 12) & to_signed(357417, 20)),
		std_logic_vector(to_signed(-1180, 12) & to_signed(356239, 20)),
		std_logic_vector(to_signed(-1183, 12) & to_signed(355057, 20)),
		std_logic_vector(to_signed(-1187, 12) & to_signed(353872, 20)),
		std_logic_vector(to_signed(-1190, 12) & to_signed(352683, 20)),
		std_logic_vector(to_signed(-1193, 12) & to_signed(351491, 20)),
		std_logic_vector(to_signed(-1197, 12) & to_signed(350296, 20)),
		std_logic_vector(to_signed(-1200, 12) & to_signed(349098, 20)),
		std_logic_vector(to_signed(-1203, 12) & to_signed(347896, 20)),
		std_logic_vector(to_signed(-1207, 12) & to_signed(346691, 20)),
		std_logic_vector(to_signed(-1210, 12) & to_signed(345483, 20)),
		std_logic_vector(to_signed(-1213, 12) & to_signed(344271, 20)),
		std_logic_vector(to_signed(-1216, 12) & to_signed(343057, 20)),
		std_logic_vector(to_signed(-1220, 12) & to_signed(341839, 20)),
		std_logic_vector(to_signed(-1223, 12) & to_signed(340618, 20)),
		std_logic_vector(to_signed(-1226, 12) & to_signed(339393, 20)),
		std_logic_vector(to_signed(-1229, 12) & to_signed(338166, 20)),
		std_logic_vector(to_signed(-1232, 12) & to_signed(336935, 20)),
		std_logic_vector(to_signed(-1236, 12) & to_signed(335701, 20)),
		std_logic_vector(to_signed(-1239, 12) & to_signed(334464, 20)),
		std_logic_vector(to_signed(-1242, 12) & to_signed(333224, 20)),
		std_logic_vector(to_signed(-1245, 12) & to_signed(331980, 20)),
		std_logic_vector(to_signed(-1248, 12) & to_signed(330734, 20)),
		std_logic_vector(to_signed(-1251, 12) & to_signed(329484, 20)),
		std_logic_vector(to_signed(-1254, 12) & to_signed(328231, 20)),
		std_logic_vector(to_signed(-1257, 12) & to_signed(326976, 20)),
		std_logic_vector(to_signed(-1260, 12) & to_signed(325717, 20)),
		std_logic_vector(to_signed(-1263, 12) & to_signed(324455, 20)),
		std_logic_vector(to_signed(-1267, 12) & to_signed(323190, 20)),
		std_logic_vector(to_signed(-1270, 12) & to_signed(321922, 20)),
		std_logic_vector(to_signed(-1273, 12) & to_signed(320651, 20)),
		std_logic_vector(to_signed(-1276, 12) & to_signed(319377, 20)),
		std_logic_vector(to_signed(-1279, 12) & to_signed(318099, 20)),
		std_logic_vector(to_signed(-1282, 12) & to_signed(316819, 20)),
		std_logic_vector(to_signed(-1285, 12) & to_signed(315536, 20)),
		std_logic_vector(to_signed(-1288, 12) & to_signed(314250, 20)),
		std_logic_vector(to_signed(-1290, 12) & to_signed(312961, 20)),
		std_logic_vector(to_signed(-1293, 12) & to_signed(311669, 20)),
		std_logic_vector(to_signed(-1296, 12) & to_signed(310374, 20)),
		std_logic_vector(to_signed(-1299, 12) & to_signed(309077, 20)),
		std_logic_vector(to_signed(-1302, 12) & to_signed(307776, 20)),
		std_logic_vector(to_signed(-1305, 12) & to_signed(306472, 20)),
		std_logic_vector(to_signed(-1308, 12) & to_signed(305166, 20)),
		std_logic_vector(to_signed(-1311, 12) & to_signed(303856, 20)),
		std_logic_vector(to_signed(-1314, 12) & to_signed(302544, 20)),
		std_logic_vector(to_signed(-1316, 12) & to_signed(301229, 20)),
		std_logic_vector(to_signed(-1319, 12) & to_signed(299911, 20)),
		std_logic_vector(to_signed(-1322, 12) & to_signed(298590, 20)),
		std_logic_vector(to_signed(-1325, 12) & to_signed(297267, 20)),
		std_logic_vector(to_signed(-1328, 12) & to_signed(295941, 20)),
		std_logic_vector(to_signed(-1331, 12) & to_signed(294611, 20)),
		std_logic_vector(to_signed(-1333, 12) & to_signed(293280, 20)),
		std_logic_vector(to_signed(-1336, 12) & to_signed(291945, 20)),
		std_logic_vector(to_signed(-1339, 12) & to_signed(290608, 20)),
		std_logic_vector(to_signed(-1342, 12) & to_signed(289267, 20)),
		std_logic_vector(to_signed(-1344, 12) & to_signed(287925, 20)),
		std_logic_vector(to_signed(-1347, 12) & to_signed(286579, 20)),
		std_logic_vector(to_signed(-1350, 12) & to_signed(285231, 20)),
		std_logic_vector(to_signed(-1352, 12) & to_signed(283880, 20)),
		std_logic_vector(to_signed(-1355, 12) & to_signed(282526, 20)),
		std_logic_vector(to_signed(-1358, 12) & to_signed(281170, 20)),
		std_logic_vector(to_signed(-1360, 12) & to_signed(279811, 20)),
		std_logic_vector(to_signed(-1363, 12) & to_signed(278449, 20)),
		std_logic_vector(to_signed(-1365, 12) & to_signed(277085, 20)),
		std_logic_vector(to_signed(-1368, 12) & to_signed(275718, 20)),
		std_logic_vector(to_signed(-1371, 12) & to_signed(274349, 20)),
		std_logic_vector(to_signed(-1373, 12) & to_signed(272977, 20)),
		std_logic_vector(to_signed(-1376, 12) & to_signed(271602, 20)),
		std_logic_vector(to_signed(-1378, 12) & to_signed(270225, 20)),
		std_logic_vector(to_signed(-1381, 12) & to_signed(268846, 20)),
		std_logic_vector(to_signed(-1383, 12) & to_signed(267464, 20)),
		std_logic_vector(to_signed(-1386, 12) & to_signed(266079, 20)),
		std_logic_vector(to_signed(-1388, 12) & to_signed(264692, 20)),
		std_logic_vector(to_signed(-1391, 12) & to_signed(263302, 20)),
		std_logic_vector(to_signed(-1393, 12) & to_signed(261910, 20)),
		std_logic_vector(to_signed(-1396, 12) & to_signed(260515, 20)),
		std_logic_vector(to_signed(-1398, 12) & to_signed(259118, 20)),
		std_logic_vector(to_signed(-1401, 12) & to_signed(257719, 20)),
		std_logic_vector(to_signed(-1403, 12) & to_signed(256317, 20)),
		std_logic_vector(to_signed(-1406, 12) & to_signed(254912, 20)),
		std_logic_vector(to_signed(-1408, 12) & to_signed(253506, 20)),
		std_logic_vector(to_signed(-1410, 12) & to_signed(252096, 20)),
		std_logic_vector(to_signed(-1413, 12) & to_signed(250685, 20)),
		std_logic_vector(to_signed(-1415, 12) & to_signed(249271, 20)),
		std_logic_vector(to_signed(-1417, 12) & to_signed(247855, 20)),
		std_logic_vector(to_signed(-1420, 12) & to_signed(246436, 20)),
		std_logic_vector(to_signed(-1422, 12) & to_signed(245015, 20)),
		std_logic_vector(to_signed(-1424, 12) & to_signed(243592, 20)),
		std_logic_vector(to_signed(-1427, 12) & to_signed(242167, 20)),
		std_logic_vector(to_signed(-1429, 12) & to_signed(240739, 20)),
		std_logic_vector(to_signed(-1431, 12) & to_signed(239309, 20)),
		std_logic_vector(to_signed(-1433, 12) & to_signed(237877, 20)),
		std_logic_vector(to_signed(-1436, 12) & to_signed(236442, 20)),
		std_logic_vector(to_signed(-1438, 12) & to_signed(235005, 20)),
		std_logic_vector(to_signed(-1440, 12) & to_signed(233566, 20)),
		std_logic_vector(to_signed(-1442, 12) & to_signed(232125, 20)),
		std_logic_vector(to_signed(-1444, 12) & to_signed(230682, 20)),
		std_logic_vector(to_signed(-1447, 12) & to_signed(229236, 20)),
		std_logic_vector(to_signed(-1449, 12) & to_signed(227789, 20)),
		std_logic_vector(to_signed(-1451, 12) & to_signed(226339, 20)),
		std_logic_vector(to_signed(-1453, 12) & to_signed(224887, 20)),
		std_logic_vector(to_signed(-1455, 12) & to_signed(223433, 20)),
		std_logic_vector(to_signed(-1457, 12) & to_signed(221977, 20)),
		std_logic_vector(to_signed(-1459, 12) & to_signed(220519, 20)),
		std_logic_vector(to_signed(-1461, 12) & to_signed(219058, 20)),
		std_logic_vector(to_signed(-1463, 12) & to_signed(217596, 20)),
		std_logic_vector(to_signed(-1465, 12) & to_signed(216131, 20)),
		std_logic_vector(to_signed(-1467, 12) & to_signed(214665, 20)),
		std_logic_vector(to_signed(-1469, 12) & to_signed(213197, 20)),
		std_logic_vector(to_signed(-1471, 12) & to_signed(211726, 20)),
		std_logic_vector(to_signed(-1473, 12) & to_signed(210254, 20)),
		std_logic_vector(to_signed(-1475, 12) & to_signed(208779, 20)),
		std_logic_vector(to_signed(-1477, 12) & to_signed(207303, 20)),
		std_logic_vector(to_signed(-1479, 12) & to_signed(205824, 20)),
		std_logic_vector(to_signed(-1481, 12) & to_signed(204344, 20)),
		std_logic_vector(to_signed(-1483, 12) & to_signed(202862, 20)),
		std_logic_vector(to_signed(-1485, 12) & to_signed(201378, 20)),
		std_logic_vector(to_signed(-1487, 12) & to_signed(199892, 20)),
		std_logic_vector(to_signed(-1489, 12) & to_signed(198404, 20)),
		std_logic_vector(to_signed(-1491, 12) & to_signed(196914, 20)),
		std_logic_vector(to_signed(-1493, 12) & to_signed(195422, 20)),
		std_logic_vector(to_signed(-1494, 12) & to_signed(193929, 20)),
		std_logic_vector(to_signed(-1496, 12) & to_signed(192433, 20)),
		std_logic_vector(to_signed(-1498, 12) & to_signed(190936, 20)),
		std_logic_vector(to_signed(-1500, 12) & to_signed(189437, 20)),
		std_logic_vector(to_signed(-1502, 12) & to_signed(187937, 20)),
		std_logic_vector(to_signed(-1503, 12) & to_signed(186434, 20)),
		std_logic_vector(to_signed(-1505, 12) & to_signed(184930, 20)),
		std_logic_vector(to_signed(-1507, 12) & to_signed(183424, 20)),
		std_logic_vector(to_signed(-1509, 12) & to_signed(181916, 20)),
		std_logic_vector(to_signed(-1510, 12) & to_signed(180407, 20)),
		std_logic_vector(to_signed(-1512, 12) & to_signed(178896, 20)),
		std_logic_vector(to_signed(-1514, 12) & to_signed(177383, 20)),
		std_logic_vector(to_signed(-1515, 12) & to_signed(175869, 20)),
		std_logic_vector(to_signed(-1517, 12) & to_signed(174352, 20)),
		std_logic_vector(to_signed(-1519, 12) & to_signed(172835, 20)),
		std_logic_vector(to_signed(-1520, 12) & to_signed(171315, 20)),
		std_logic_vector(to_signed(-1522, 12) & to_signed(169794, 20)),
		std_logic_vector(to_signed(-1523, 12) & to_signed(168272, 20)),
		std_logic_vector(to_signed(-1525, 12) & to_signed(166748, 20)),
		std_logic_vector(to_signed(-1527, 12) & to_signed(165222, 20)),
		std_logic_vector(to_signed(-1528, 12) & to_signed(163694, 20)),
		std_logic_vector(to_signed(-1530, 12) & to_signed(162166, 20)),
		std_logic_vector(to_signed(-1531, 12) & to_signed(160635, 20)),
		std_logic_vector(to_signed(-1533, 12) & to_signed(159103, 20)),
		std_logic_vector(to_signed(-1534, 12) & to_signed(157570, 20)),
		std_logic_vector(to_signed(-1536, 12) & to_signed(156035, 20)),
		std_logic_vector(to_signed(-1537, 12) & to_signed(154499, 20)),
		std_logic_vector(to_signed(-1539, 12) & to_signed(152961, 20)),
		std_logic_vector(to_signed(-1540, 12) & to_signed(151422, 20)),
		std_logic_vector(to_signed(-1541, 12) & to_signed(149881, 20)),
		std_logic_vector(to_signed(-1543, 12) & to_signed(148339, 20)),
		std_logic_vector(to_signed(-1544, 12) & to_signed(146796, 20)),
		std_logic_vector(to_signed(-1546, 12) & to_signed(145251, 20)),
		std_logic_vector(to_signed(-1547, 12) & to_signed(143705, 20)),
		std_logic_vector(to_signed(-1548, 12) & to_signed(142157, 20)),
		std_logic_vector(to_signed(-1550, 12) & to_signed(140608, 20)),
		std_logic_vector(to_signed(-1551, 12) & to_signed(139058, 20)),
		std_logic_vector(to_signed(-1552, 12) & to_signed(137506, 20)),
		std_logic_vector(to_signed(-1553, 12) & to_signed(135954, 20)),
		std_logic_vector(to_signed(-1555, 12) & to_signed(134400, 20)),
		std_logic_vector(to_signed(-1556, 12) & to_signed(132844, 20)),
		std_logic_vector(to_signed(-1557, 12) & to_signed(131288, 20)),
		std_logic_vector(to_signed(-1558, 12) & to_signed(129730, 20)),
		std_logic_vector(to_signed(-1560, 12) & to_signed(128171, 20)),
		std_logic_vector(to_signed(-1561, 12) & to_signed(126610, 20)),
		std_logic_vector(to_signed(-1562, 12) & to_signed(125049, 20)),
		std_logic_vector(to_signed(-1563, 12) & to_signed(123486, 20)),
		std_logic_vector(to_signed(-1564, 12) & to_signed(121922, 20)),
		std_logic_vector(to_signed(-1566, 12) & to_signed(120357, 20)),
		std_logic_vector(to_signed(-1567, 12) & to_signed(118791, 20)),
		std_logic_vector(to_signed(-1568, 12) & to_signed(117224, 20)),
		std_logic_vector(to_signed(-1569, 12) & to_signed(115656, 20)),
		std_logic_vector(to_signed(-1570, 12) & to_signed(114086, 20)),
		std_logic_vector(to_signed(-1571, 12) & to_signed(112516, 20)),
		std_logic_vector(to_signed(-1572, 12) & to_signed(110944, 20)),
		std_logic_vector(to_signed(-1573, 12) & to_signed(109372, 20)),
		std_logic_vector(to_signed(-1574, 12) & to_signed(107798, 20)),
		std_logic_vector(to_signed(-1575, 12) & to_signed(106224, 20)),
		std_logic_vector(to_signed(-1576, 12) & to_signed(104648, 20)),
		std_logic_vector(to_signed(-1577, 12) & to_signed(103071, 20)),
		std_logic_vector(to_signed(-1578, 12) & to_signed(101494, 20)),
		std_logic_vector(to_signed(-1579, 12) & to_signed(99915, 20)),
		std_logic_vector(to_signed(-1580, 12) & to_signed(98336, 20)),
		std_logic_vector(to_signed(-1581, 12) & to_signed(96755, 20)),
		std_logic_vector(to_signed(-1582, 12) & to_signed(95174, 20)),
		std_logic_vector(to_signed(-1583, 12) & to_signed(93592, 20)),
		std_logic_vector(to_signed(-1584, 12) & to_signed(92009, 20)),
		std_logic_vector(to_signed(-1584, 12) & to_signed(90425, 20)),
		std_logic_vector(to_signed(-1585, 12) & to_signed(88840, 20)),
		std_logic_vector(to_signed(-1586, 12) & to_signed(87254, 20)),
		std_logic_vector(to_signed(-1587, 12) & to_signed(85668, 20)),
		std_logic_vector(to_signed(-1588, 12) & to_signed(84081, 20)),
		std_logic_vector(to_signed(-1588, 12) & to_signed(82493, 20)),
		std_logic_vector(to_signed(-1589, 12) & to_signed(80904, 20)),
		std_logic_vector(to_signed(-1590, 12) & to_signed(79314, 20)),
		std_logic_vector(to_signed(-1591, 12) & to_signed(77724, 20)),
		std_logic_vector(to_signed(-1591, 12) & to_signed(76133, 20)),
		std_logic_vector(to_signed(-1592, 12) & to_signed(74541, 20)),
		std_logic_vector(to_signed(-1593, 12) & to_signed(72949, 20)),
		std_logic_vector(to_signed(-1594, 12) & to_signed(71355, 20)),
		std_logic_vector(to_signed(-1594, 12) & to_signed(69762, 20)),
		std_logic_vector(to_signed(-1595, 12) & to_signed(68167, 20)),
		std_logic_vector(to_signed(-1595, 12) & to_signed(66572, 20)),
		std_logic_vector(to_signed(-1596, 12) & to_signed(64976, 20)),
		std_logic_vector(to_signed(-1597, 12) & to_signed(63380, 20)),
		std_logic_vector(to_signed(-1597, 12) & to_signed(61783, 20)),
		std_logic_vector(to_signed(-1598, 12) & to_signed(60185, 20)),
		std_logic_vector(to_signed(-1598, 12) & to_signed(58587, 20)),
		std_logic_vector(to_signed(-1599, 12) & to_signed(56988, 20)),
		std_logic_vector(to_signed(-1599, 12) & to_signed(55389, 20)),
		std_logic_vector(to_signed(-1600, 12) & to_signed(53789, 20)),
		std_logic_vector(to_signed(-1600, 12) & to_signed(52189, 20)),
		std_logic_vector(to_signed(-1601, 12) & to_signed(50588, 20)),
		std_logic_vector(to_signed(-1601, 12) & to_signed(48987, 20)),
		std_logic_vector(to_signed(-1602, 12) & to_signed(47386, 20)),
		std_logic_vector(to_signed(-1602, 12) & to_signed(45783, 20)),
		std_logic_vector(to_signed(-1603, 12) & to_signed(44181, 20)),
		std_logic_vector(to_signed(-1603, 12) & to_signed(42578, 20)),
		std_logic_vector(to_signed(-1604, 12) & to_signed(40974, 20)),
		std_logic_vector(to_signed(-1604, 12) & to_signed(39371, 20)),
		std_logic_vector(to_signed(-1604, 12) & to_signed(37767, 20)),
		std_logic_vector(to_signed(-1605, 12) & to_signed(36162, 20)),
		std_logic_vector(to_signed(-1605, 12) & to_signed(34557, 20)),
		std_logic_vector(to_signed(-1605, 12) & to_signed(32952, 20)),
		std_logic_vector(to_signed(-1606, 12) & to_signed(31347, 20)),
		std_logic_vector(to_signed(-1606, 12) & to_signed(29741, 20)),
		std_logic_vector(to_signed(-1606, 12) & to_signed(28135, 20)),
		std_logic_vector(to_signed(-1606, 12) & to_signed(26529, 20)),
		std_logic_vector(to_signed(-1607, 12) & to_signed(24922, 20)),
		std_logic_vector(to_signed(-1607, 12) & to_signed(23315, 20)),
		std_logic_vector(to_signed(-1607, 12) & to_signed(21708, 20)),
		std_logic_vector(to_signed(-1607, 12) & to_signed(20101, 20)),
		std_logic_vector(to_signed(-1607, 12) & to_signed(18494, 20)),
		std_logic_vector(to_signed(-1608, 12) & to_signed(16886, 20)),
		std_logic_vector(to_signed(-1608, 12) & to_signed(15278, 20)),
		std_logic_vector(to_signed(-1608, 12) & to_signed(13671, 20)),
		std_logic_vector(to_signed(-1608, 12) & to_signed(12063, 20)),
		std_logic_vector(to_signed(-1608, 12) & to_signed(10454, 20)),
		std_logic_vector(to_signed(-1608, 12) & to_signed(8846, 20)),
		std_logic_vector(to_signed(-1608, 12) & to_signed(7238, 20)),
		std_logic_vector(to_signed(-1608, 12) & to_signed(5630, 20)),
		std_logic_vector(to_signed(-1608, 12) & to_signed(4021, 20)),
		std_logic_vector(to_signed(-1608, 12) & to_signed(2413, 20)),
		std_logic_vector(to_signed(-1608, 12) & to_signed(804, 20)),
		std_logic_vector(to_signed(-1608, 12) & to_signed(-804, 20)),
		std_logic_vector(to_signed(-1608, 12) & to_signed(-2413, 20)),
		std_logic_vector(to_signed(-1608, 12) & to_signed(-4021, 20)),
		std_logic_vector(to_signed(-1608, 12) & to_signed(-5630, 20)),
		std_logic_vector(to_signed(-1608, 12) & to_signed(-7238, 20)),
		std_logic_vector(to_signed(-1608, 12) & to_signed(-8846, 20)),
		std_logic_vector(to_signed(-1608, 12) & to_signed(-10454, 20)),
		std_logic_vector(to_signed(-1608, 12) & to_signed(-12063, 20)),
		std_logic_vector(to_signed(-1608, 12) & to_signed(-13671, 20)),
		std_logic_vector(to_signed(-1608, 12) & to_signed(-15278, 20)),
		std_logic_vector(to_signed(-1608, 12) & to_signed(-16886, 20)),
		std_logic_vector(to_signed(-1607, 12) & to_signed(-18494, 20)),
		std_logic_vector(to_signed(-1607, 12) & to_signed(-20101, 20)),
		std_logic_vector(to_signed(-1607, 12) & to_signed(-21708, 20)),
		std_logic_vector(to_signed(-1607, 12) & to_signed(-23315, 20)),
		std_logic_vector(to_signed(-1607, 12) & to_signed(-24922, 20)),
		std_logic_vector(to_signed(-1606, 12) & to_signed(-26529, 20)),
		std_logic_vector(to_signed(-1606, 12) & to_signed(-28135, 20)),
		std_logic_vector(to_signed(-1606, 12) & to_signed(-29741, 20)),
		std_logic_vector(to_signed(-1606, 12) & to_signed(-31347, 20)),
		std_logic_vector(to_signed(-1605, 12) & to_signed(-32952, 20)),
		std_logic_vector(to_signed(-1605, 12) & to_signed(-34557, 20)),
		std_logic_vector(to_signed(-1605, 12) & to_signed(-36162, 20)),
		std_logic_vector(to_signed(-1604, 12) & to_signed(-37767, 20)),
		std_logic_vector(to_signed(-1604, 12) & to_signed(-39371, 20)),
		std_logic_vector(to_signed(-1604, 12) & to_signed(-40974, 20)),
		std_logic_vector(to_signed(-1603, 12) & to_signed(-42578, 20)),
		std_logic_vector(to_signed(-1603, 12) & to_signed(-44181, 20)),
		std_logic_vector(to_signed(-1602, 12) & to_signed(-45783, 20)),
		std_logic_vector(to_signed(-1602, 12) & to_signed(-47386, 20)),
		std_logic_vector(to_signed(-1601, 12) & to_signed(-48987, 20)),
		std_logic_vector(to_signed(-1601, 12) & to_signed(-50588, 20)),
		std_logic_vector(to_signed(-1600, 12) & to_signed(-52189, 20)),
		std_logic_vector(to_signed(-1600, 12) & to_signed(-53789, 20)),
		std_logic_vector(to_signed(-1599, 12) & to_signed(-55389, 20)),
		std_logic_vector(to_signed(-1599, 12) & to_signed(-56988, 20)),
		std_logic_vector(to_signed(-1598, 12) & to_signed(-58587, 20)),
		std_logic_vector(to_signed(-1598, 12) & to_signed(-60185, 20)),
		std_logic_vector(to_signed(-1597, 12) & to_signed(-61783, 20)),
		std_logic_vector(to_signed(-1597, 12) & to_signed(-63380, 20)),
		std_logic_vector(to_signed(-1596, 12) & to_signed(-64976, 20)),
		std_logic_vector(to_signed(-1595, 12) & to_signed(-66572, 20)),
		std_logic_vector(to_signed(-1595, 12) & to_signed(-68167, 20)),
		std_logic_vector(to_signed(-1594, 12) & to_signed(-69762, 20)),
		std_logic_vector(to_signed(-1594, 12) & to_signed(-71355, 20)),
		std_logic_vector(to_signed(-1593, 12) & to_signed(-72949, 20)),
		std_logic_vector(to_signed(-1592, 12) & to_signed(-74541, 20)),
		std_logic_vector(to_signed(-1591, 12) & to_signed(-76133, 20)),
		std_logic_vector(to_signed(-1591, 12) & to_signed(-77724, 20)),
		std_logic_vector(to_signed(-1590, 12) & to_signed(-79314, 20)),
		std_logic_vector(to_signed(-1589, 12) & to_signed(-80904, 20)),
		std_logic_vector(to_signed(-1588, 12) & to_signed(-82493, 20)),
		std_logic_vector(to_signed(-1588, 12) & to_signed(-84081, 20)),
		std_logic_vector(to_signed(-1587, 12) & to_signed(-85668, 20)),
		std_logic_vector(to_signed(-1586, 12) & to_signed(-87254, 20)),
		std_logic_vector(to_signed(-1585, 12) & to_signed(-88840, 20)),
		std_logic_vector(to_signed(-1584, 12) & to_signed(-90425, 20)),
		std_logic_vector(to_signed(-1584, 12) & to_signed(-92009, 20)),
		std_logic_vector(to_signed(-1583, 12) & to_signed(-93592, 20)),
		std_logic_vector(to_signed(-1582, 12) & to_signed(-95174, 20)),
		std_logic_vector(to_signed(-1581, 12) & to_signed(-96755, 20)),
		std_logic_vector(to_signed(-1580, 12) & to_signed(-98336, 20)),
		std_logic_vector(to_signed(-1579, 12) & to_signed(-99915, 20)),
		std_logic_vector(to_signed(-1578, 12) & to_signed(-101494, 20)),
		std_logic_vector(to_signed(-1577, 12) & to_signed(-103071, 20)),
		std_logic_vector(to_signed(-1576, 12) & to_signed(-104648, 20)),
		std_logic_vector(to_signed(-1575, 12) & to_signed(-106224, 20)),
		std_logic_vector(to_signed(-1574, 12) & to_signed(-107798, 20)),
		std_logic_vector(to_signed(-1573, 12) & to_signed(-109372, 20)),
		std_logic_vector(to_signed(-1572, 12) & to_signed(-110944, 20)),
		std_logic_vector(to_signed(-1571, 12) & to_signed(-112516, 20)),
		std_logic_vector(to_signed(-1570, 12) & to_signed(-114086, 20)),
		std_logic_vector(to_signed(-1569, 12) & to_signed(-115656, 20)),
		std_logic_vector(to_signed(-1568, 12) & to_signed(-117224, 20)),
		std_logic_vector(to_signed(-1567, 12) & to_signed(-118791, 20)),
		std_logic_vector(to_signed(-1566, 12) & to_signed(-120357, 20)),
		std_logic_vector(to_signed(-1564, 12) & to_signed(-121922, 20)),
		std_logic_vector(to_signed(-1563, 12) & to_signed(-123486, 20)),
		std_logic_vector(to_signed(-1562, 12) & to_signed(-125049, 20)),
		std_logic_vector(to_signed(-1561, 12) & to_signed(-126610, 20)),
		std_logic_vector(to_signed(-1560, 12) & to_signed(-128171, 20)),
		std_logic_vector(to_signed(-1558, 12) & to_signed(-129730, 20)),
		std_logic_vector(to_signed(-1557, 12) & to_signed(-131288, 20)),
		std_logic_vector(to_signed(-1556, 12) & to_signed(-132844, 20)),
		std_logic_vector(to_signed(-1555, 12) & to_signed(-134400, 20)),
		std_logic_vector(to_signed(-1553, 12) & to_signed(-135954, 20)),
		std_logic_vector(to_signed(-1552, 12) & to_signed(-137506, 20)),
		std_logic_vector(to_signed(-1551, 12) & to_signed(-139058, 20)),
		std_logic_vector(to_signed(-1550, 12) & to_signed(-140608, 20)),
		std_logic_vector(to_signed(-1548, 12) & to_signed(-142157, 20)),
		std_logic_vector(to_signed(-1547, 12) & to_signed(-143705, 20)),
		std_logic_vector(to_signed(-1546, 12) & to_signed(-145251, 20)),
		std_logic_vector(to_signed(-1544, 12) & to_signed(-146796, 20)),
		std_logic_vector(to_signed(-1543, 12) & to_signed(-148339, 20)),
		std_logic_vector(to_signed(-1541, 12) & to_signed(-149881, 20)),
		std_logic_vector(to_signed(-1540, 12) & to_signed(-151422, 20)),
		std_logic_vector(to_signed(-1539, 12) & to_signed(-152961, 20)),
		std_logic_vector(to_signed(-1537, 12) & to_signed(-154499, 20)),
		std_logic_vector(to_signed(-1536, 12) & to_signed(-156035, 20)),
		std_logic_vector(to_signed(-1534, 12) & to_signed(-157570, 20)),
		std_logic_vector(to_signed(-1533, 12) & to_signed(-159103, 20)),
		std_logic_vector(to_signed(-1531, 12) & to_signed(-160635, 20)),
		std_logic_vector(to_signed(-1530, 12) & to_signed(-162166, 20)),
		std_logic_vector(to_signed(-1528, 12) & to_signed(-163694, 20)),
		std_logic_vector(to_signed(-1527, 12) & to_signed(-165222, 20)),
		std_logic_vector(to_signed(-1525, 12) & to_signed(-166748, 20)),
		std_logic_vector(to_signed(-1523, 12) & to_signed(-168272, 20)),
		std_logic_vector(to_signed(-1522, 12) & to_signed(-169794, 20)),
		std_logic_vector(to_signed(-1520, 12) & to_signed(-171315, 20)),
		std_logic_vector(to_signed(-1519, 12) & to_signed(-172835, 20)),
		std_logic_vector(to_signed(-1517, 12) & to_signed(-174352, 20)),
		std_logic_vector(to_signed(-1515, 12) & to_signed(-175869, 20)),
		std_logic_vector(to_signed(-1514, 12) & to_signed(-177383, 20)),
		std_logic_vector(to_signed(-1512, 12) & to_signed(-178896, 20)),
		std_logic_vector(to_signed(-1510, 12) & to_signed(-180407, 20)),
		std_logic_vector(to_signed(-1509, 12) & to_signed(-181916, 20)),
		std_logic_vector(to_signed(-1507, 12) & to_signed(-183424, 20)),
		std_logic_vector(to_signed(-1505, 12) & to_signed(-184930, 20)),
		std_logic_vector(to_signed(-1503, 12) & to_signed(-186434, 20)),
		std_logic_vector(to_signed(-1502, 12) & to_signed(-187937, 20)),
		std_logic_vector(to_signed(-1500, 12) & to_signed(-189437, 20)),
		std_logic_vector(to_signed(-1498, 12) & to_signed(-190936, 20)),
		std_logic_vector(to_signed(-1496, 12) & to_signed(-192433, 20)),
		std_logic_vector(to_signed(-1494, 12) & to_signed(-193929, 20)),
		std_logic_vector(to_signed(-1493, 12) & to_signed(-195422, 20)),
		std_logic_vector(to_signed(-1491, 12) & to_signed(-196914, 20)),
		std_logic_vector(to_signed(-1489, 12) & to_signed(-198404, 20)),
		std_logic_vector(to_signed(-1487, 12) & to_signed(-199892, 20)),
		std_logic_vector(to_signed(-1485, 12) & to_signed(-201378, 20)),
		std_logic_vector(to_signed(-1483, 12) & to_signed(-202862, 20)),
		std_logic_vector(to_signed(-1481, 12) & to_signed(-204344, 20)),
		std_logic_vector(to_signed(-1479, 12) & to_signed(-205824, 20)),
		std_logic_vector(to_signed(-1477, 12) & to_signed(-207303, 20)),
		std_logic_vector(to_signed(-1475, 12) & to_signed(-208779, 20)),
		std_logic_vector(to_signed(-1473, 12) & to_signed(-210254, 20)),
		std_logic_vector(to_signed(-1471, 12) & to_signed(-211726, 20)),
		std_logic_vector(to_signed(-1469, 12) & to_signed(-213197, 20)),
		std_logic_vector(to_signed(-1467, 12) & to_signed(-214665, 20)),
		std_logic_vector(to_signed(-1465, 12) & to_signed(-216131, 20)),
		std_logic_vector(to_signed(-1463, 12) & to_signed(-217596, 20)),
		std_logic_vector(to_signed(-1461, 12) & to_signed(-219058, 20)),
		std_logic_vector(to_signed(-1459, 12) & to_signed(-220519, 20)),
		std_logic_vector(to_signed(-1457, 12) & to_signed(-221977, 20)),
		std_logic_vector(to_signed(-1455, 12) & to_signed(-223433, 20)),
		std_logic_vector(to_signed(-1453, 12) & to_signed(-224887, 20)),
		std_logic_vector(to_signed(-1451, 12) & to_signed(-226339, 20)),
		std_logic_vector(to_signed(-1449, 12) & to_signed(-227789, 20)),
		std_logic_vector(to_signed(-1447, 12) & to_signed(-229236, 20)),
		std_logic_vector(to_signed(-1444, 12) & to_signed(-230682, 20)),
		std_logic_vector(to_signed(-1442, 12) & to_signed(-232125, 20)),
		std_logic_vector(to_signed(-1440, 12) & to_signed(-233566, 20)),
		std_logic_vector(to_signed(-1438, 12) & to_signed(-235005, 20)),
		std_logic_vector(to_signed(-1436, 12) & to_signed(-236442, 20)),
		std_logic_vector(to_signed(-1433, 12) & to_signed(-237877, 20)),
		std_logic_vector(to_signed(-1431, 12) & to_signed(-239309, 20)),
		std_logic_vector(to_signed(-1429, 12) & to_signed(-240739, 20)),
		std_logic_vector(to_signed(-1427, 12) & to_signed(-242167, 20)),
		std_logic_vector(to_signed(-1424, 12) & to_signed(-243592, 20)),
		std_logic_vector(to_signed(-1422, 12) & to_signed(-245015, 20)),
		std_logic_vector(to_signed(-1420, 12) & to_signed(-246436, 20)),
		std_logic_vector(to_signed(-1417, 12) & to_signed(-247855, 20)),
		std_logic_vector(to_signed(-1415, 12) & to_signed(-249271, 20)),
		std_logic_vector(to_signed(-1413, 12) & to_signed(-250685, 20)),
		std_logic_vector(to_signed(-1410, 12) & to_signed(-252096, 20)),
		std_logic_vector(to_signed(-1408, 12) & to_signed(-253506, 20)),
		std_logic_vector(to_signed(-1406, 12) & to_signed(-254912, 20)),
		std_logic_vector(to_signed(-1403, 12) & to_signed(-256317, 20)),
		std_logic_vector(to_signed(-1401, 12) & to_signed(-257719, 20)),
		std_logic_vector(to_signed(-1398, 12) & to_signed(-259118, 20)),
		std_logic_vector(to_signed(-1396, 12) & to_signed(-260515, 20)),
		std_logic_vector(to_signed(-1393, 12) & to_signed(-261910, 20)),
		std_logic_vector(to_signed(-1391, 12) & to_signed(-263302, 20)),
		std_logic_vector(to_signed(-1388, 12) & to_signed(-264692, 20)),
		std_logic_vector(to_signed(-1386, 12) & to_signed(-266079, 20)),
		std_logic_vector(to_signed(-1383, 12) & to_signed(-267464, 20)),
		std_logic_vector(to_signed(-1381, 12) & to_signed(-268846, 20)),
		std_logic_vector(to_signed(-1378, 12) & to_signed(-270225, 20)),
		std_logic_vector(to_signed(-1376, 12) & to_signed(-271602, 20)),
		std_logic_vector(to_signed(-1373, 12) & to_signed(-272977, 20)),
		std_logic_vector(to_signed(-1371, 12) & to_signed(-274349, 20)),
		std_logic_vector(to_signed(-1368, 12) & to_signed(-275718, 20)),
		std_logic_vector(to_signed(-1365, 12) & to_signed(-277085, 20)),
		std_logic_vector(to_signed(-1363, 12) & to_signed(-278449, 20)),
		std_logic_vector(to_signed(-1360, 12) & to_signed(-279811, 20)),
		std_logic_vector(to_signed(-1358, 12) & to_signed(-281170, 20)),
		std_logic_vector(to_signed(-1355, 12) & to_signed(-282526, 20)),
		std_logic_vector(to_signed(-1352, 12) & to_signed(-283880, 20)),
		std_logic_vector(to_signed(-1350, 12) & to_signed(-285231, 20)),
		std_logic_vector(to_signed(-1347, 12) & to_signed(-286579, 20)),
		std_logic_vector(to_signed(-1344, 12) & to_signed(-287925, 20)),
		std_logic_vector(to_signed(-1342, 12) & to_signed(-289267, 20)),
		std_logic_vector(to_signed(-1339, 12) & to_signed(-290608, 20)),
		std_logic_vector(to_signed(-1336, 12) & to_signed(-291945, 20)),
		std_logic_vector(to_signed(-1333, 12) & to_signed(-293280, 20)),
		std_logic_vector(to_signed(-1331, 12) & to_signed(-294611, 20)),
		std_logic_vector(to_signed(-1328, 12) & to_signed(-295941, 20)),
		std_logic_vector(to_signed(-1325, 12) & to_signed(-297267, 20)),
		std_logic_vector(to_signed(-1322, 12) & to_signed(-298590, 20)),
		std_logic_vector(to_signed(-1319, 12) & to_signed(-299911, 20)),
		std_logic_vector(to_signed(-1316, 12) & to_signed(-301229, 20)),
		std_logic_vector(to_signed(-1314, 12) & to_signed(-302544, 20)),
		std_logic_vector(to_signed(-1311, 12) & to_signed(-303856, 20)),
		std_logic_vector(to_signed(-1308, 12) & to_signed(-305166, 20)),
		std_logic_vector(to_signed(-1305, 12) & to_signed(-306472, 20)),
		std_logic_vector(to_signed(-1302, 12) & to_signed(-307776, 20)),
		std_logic_vector(to_signed(-1299, 12) & to_signed(-309077, 20)),
		std_logic_vector(to_signed(-1296, 12) & to_signed(-310374, 20)),
		std_logic_vector(to_signed(-1293, 12) & to_signed(-311669, 20)),
		std_logic_vector(to_signed(-1290, 12) & to_signed(-312961, 20)),
		std_logic_vector(to_signed(-1288, 12) & to_signed(-314250, 20)),
		std_logic_vector(to_signed(-1285, 12) & to_signed(-315536, 20)),
		std_logic_vector(to_signed(-1282, 12) & to_signed(-316819, 20)),
		std_logic_vector(to_signed(-1279, 12) & to_signed(-318099, 20)),
		std_logic_vector(to_signed(-1276, 12) & to_signed(-319377, 20)),
		std_logic_vector(to_signed(-1273, 12) & to_signed(-320651, 20)),
		std_logic_vector(to_signed(-1270, 12) & to_signed(-321922, 20)),
		std_logic_vector(to_signed(-1267, 12) & to_signed(-323190, 20)),
		std_logic_vector(to_signed(-1263, 12) & to_signed(-324455, 20)),
		std_logic_vector(to_signed(-1260, 12) & to_signed(-325717, 20)),
		std_logic_vector(to_signed(-1257, 12) & to_signed(-326976, 20)),
		std_logic_vector(to_signed(-1254, 12) & to_signed(-328231, 20)),
		std_logic_vector(to_signed(-1251, 12) & to_signed(-329484, 20)),
		std_logic_vector(to_signed(-1248, 12) & to_signed(-330734, 20)),
		std_logic_vector(to_signed(-1245, 12) & to_signed(-331980, 20)),
		std_logic_vector(to_signed(-1242, 12) & to_signed(-333224, 20)),
		std_logic_vector(to_signed(-1239, 12) & to_signed(-334464, 20)),
		std_logic_vector(to_signed(-1236, 12) & to_signed(-335701, 20)),
		std_logic_vector(to_signed(-1232, 12) & to_signed(-336935, 20)),
		std_logic_vector(to_signed(-1229, 12) & to_signed(-338166, 20)),
		std_logic_vector(to_signed(-1226, 12) & to_signed(-339393, 20)),
		std_logic_vector(to_signed(-1223, 12) & to_signed(-340618, 20)),
		std_logic_vector(to_signed(-1220, 12) & to_signed(-341839, 20)),
		std_logic_vector(to_signed(-1216, 12) & to_signed(-343057, 20)),
		std_logic_vector(to_signed(-1213, 12) & to_signed(-344271, 20)),
		std_logic_vector(to_signed(-1210, 12) & to_signed(-345483, 20)),
		std_logic_vector(to_signed(-1207, 12) & to_signed(-346691, 20)),
		std_logic_vector(to_signed(-1203, 12) & to_signed(-347896, 20)),
		std_logic_vector(to_signed(-1200, 12) & to_signed(-349098, 20)),
		std_logic_vector(to_signed(-1197, 12) & to_signed(-350296, 20)),
		std_logic_vector(to_signed(-1193, 12) & to_signed(-351491, 20)),
		std_logic_vector(to_signed(-1190, 12) & to_signed(-352683, 20)),
		std_logic_vector(to_signed(-1187, 12) & to_signed(-353872, 20)),
		std_logic_vector(to_signed(-1183, 12) & to_signed(-355057, 20)),
		std_logic_vector(to_signed(-1180, 12) & to_signed(-356239, 20)),
		std_logic_vector(to_signed(-1177, 12) & to_signed(-357417, 20)),
		std_logic_vector(to_signed(-1173, 12) & to_signed(-358592, 20)),
		std_logic_vector(to_signed(-1170, 12) & to_signed(-359764, 20)),
		std_logic_vector(to_signed(-1167, 12) & to_signed(-360932, 20)),
		std_logic_vector(to_signed(-1163, 12) & to_signed(-362097, 20)),
		std_logic_vector(to_signed(-1160, 12) & to_signed(-363259, 20)),
		std_logic_vector(to_signed(-1156, 12) & to_signed(-364417, 20)),
		std_logic_vector(to_signed(-1153, 12) & to_signed(-365571, 20)),
		std_logic_vector(to_signed(-1150, 12) & to_signed(-366723, 20)),
		std_logic_vector(to_signed(-1146, 12) & to_signed(-367870, 20)),
		std_logic_vector(to_signed(-1143, 12) & to_signed(-369015, 20)),
		std_logic_vector(to_signed(-1139, 12) & to_signed(-370156, 20)),
		std_logic_vector(to_signed(-1136, 12) & to_signed(-371293, 20)),
		std_logic_vector(to_signed(-1132, 12) & to_signed(-372427, 20)),
		std_logic_vector(to_signed(-1129, 12) & to_signed(-373557, 20)),
		std_logic_vector(to_signed(-1125, 12) & to_signed(-374684, 20)),
		std_logic_vector(to_signed(-1122, 12) & to_signed(-375807, 20)),
		std_logic_vector(to_signed(-1118, 12) & to_signed(-376927, 20)),
		std_logic_vector(to_signed(-1114, 12) & to_signed(-378043, 20)),
		std_logic_vector(to_signed(-1111, 12) & to_signed(-379156, 20)),
		std_logic_vector(to_signed(-1107, 12) & to_signed(-380265, 20)),
		std_logic_vector(to_signed(-1104, 12) & to_signed(-381371, 20)),
		std_logic_vector(to_signed(-1100, 12) & to_signed(-382473, 20)),
		std_logic_vector(to_signed(-1097, 12) & to_signed(-383571, 20)),
		std_logic_vector(to_signed(-1093, 12) & to_signed(-384666, 20)),
		std_logic_vector(to_signed(-1089, 12) & to_signed(-385757, 20)),
		std_logic_vector(to_signed(-1086, 12) & to_signed(-386844, 20)),
		std_logic_vector(to_signed(-1082, 12) & to_signed(-387928, 20)),
		std_logic_vector(to_signed(-1078, 12) & to_signed(-389008, 20)),
		std_logic_vector(to_signed(-1075, 12) & to_signed(-390085, 20)),
		std_logic_vector(to_signed(-1071, 12) & to_signed(-391158, 20)),
		std_logic_vector(to_signed(-1067, 12) & to_signed(-392227, 20)),
		std_logic_vector(to_signed(-1064, 12) & to_signed(-393293, 20)),
		std_logic_vector(to_signed(-1060, 12) & to_signed(-394354, 20)),
		std_logic_vector(to_signed(-1056, 12) & to_signed(-395412, 20)),
		std_logic_vector(to_signed(-1052, 12) & to_signed(-396467, 20)),
		std_logic_vector(to_signed(-1049, 12) & to_signed(-397517, 20)),
		std_logic_vector(to_signed(-1045, 12) & to_signed(-398564, 20)),
		std_logic_vector(to_signed(-1041, 12) & to_signed(-399607, 20)),
		std_logic_vector(to_signed(-1037, 12) & to_signed(-400647, 20)),
		std_logic_vector(to_signed(-1034, 12) & to_signed(-401682, 20)),
		std_logic_vector(to_signed(-1030, 12) & to_signed(-402714, 20)),
		std_logic_vector(to_signed(-1026, 12) & to_signed(-403742, 20)),
		std_logic_vector(to_signed(-1022, 12) & to_signed(-404766, 20)),
		std_logic_vector(to_signed(-1019, 12) & to_signed(-405787, 20)),
		std_logic_vector(to_signed(-1015, 12) & to_signed(-406803, 20)),
		std_logic_vector(to_signed(-1011, 12) & to_signed(-407816, 20)),
		std_logic_vector(to_signed(-1007, 12) & to_signed(-408825, 20)),
		std_logic_vector(to_signed(-1003, 12) & to_signed(-409830, 20)),
		std_logic_vector(to_signed(-999, 12) & to_signed(-410831, 20)),
		std_logic_vector(to_signed(-995, 12) & to_signed(-411829, 20)),
		std_logic_vector(to_signed(-992, 12) & to_signed(-412822, 20)),
		std_logic_vector(to_signed(-988, 12) & to_signed(-413812, 20)),
		std_logic_vector(to_signed(-984, 12) & to_signed(-414797, 20)),
		std_logic_vector(to_signed(-980, 12) & to_signed(-415779, 20)),
		std_logic_vector(to_signed(-976, 12) & to_signed(-416757, 20)),
		std_logic_vector(to_signed(-972, 12) & to_signed(-417731, 20)),
		std_logic_vector(to_signed(-968, 12) & to_signed(-418701, 20)),
		std_logic_vector(to_signed(-964, 12) & to_signed(-419667, 20)),
		std_logic_vector(to_signed(-960, 12) & to_signed(-420629, 20)),
		std_logic_vector(to_signed(-956, 12) & to_signed(-421587, 20)),
		std_logic_vector(to_signed(-952, 12) & to_signed(-422542, 20)),
		std_logic_vector(to_signed(-948, 12) & to_signed(-423492, 20)),
		std_logic_vector(to_signed(-944, 12) & to_signed(-424438, 20)),
		std_logic_vector(to_signed(-940, 12) & to_signed(-425380, 20)),
		std_logic_vector(to_signed(-936, 12) & to_signed(-426319, 20)),
		std_logic_vector(to_signed(-932, 12) & to_signed(-427253, 20)),
		std_logic_vector(to_signed(-928, 12) & to_signed(-428183, 20)),
		std_logic_vector(to_signed(-924, 12) & to_signed(-429109, 20)),
		std_logic_vector(to_signed(-920, 12) & to_signed(-430031, 20)),
		std_logic_vector(to_signed(-916, 12) & to_signed(-430949, 20)),
		std_logic_vector(to_signed(-912, 12) & to_signed(-431863, 20)),
		std_logic_vector(to_signed(-908, 12) & to_signed(-432773, 20)),
		std_logic_vector(to_signed(-904, 12) & to_signed(-433679, 20)),
		std_logic_vector(to_signed(-900, 12) & to_signed(-434581, 20)),
		std_logic_vector(to_signed(-896, 12) & to_signed(-435479, 20)),
		std_logic_vector(to_signed(-892, 12) & to_signed(-436373, 20)),
		std_logic_vector(to_signed(-887, 12) & to_signed(-437262, 20)),
		std_logic_vector(to_signed(-883, 12) & to_signed(-438147, 20)),
		std_logic_vector(to_signed(-879, 12) & to_signed(-439029, 20)),
		std_logic_vector(to_signed(-875, 12) & to_signed(-439906, 20)),
		std_logic_vector(to_signed(-871, 12) & to_signed(-440779, 20)),
		std_logic_vector(to_signed(-867, 12) & to_signed(-441648, 20)),
		std_logic_vector(to_signed(-863, 12) & to_signed(-442512, 20)),
		std_logic_vector(to_signed(-858, 12) & to_signed(-443373, 20)),
		std_logic_vector(to_signed(-854, 12) & to_signed(-444229, 20)),
		std_logic_vector(to_signed(-850, 12) & to_signed(-445081, 20)),
		std_logic_vector(to_signed(-846, 12) & to_signed(-445929, 20)),
		std_logic_vector(to_signed(-842, 12) & to_signed(-446773, 20)),
		std_logic_vector(to_signed(-837, 12) & to_signed(-447613, 20)),
		std_logic_vector(to_signed(-833, 12) & to_signed(-448448, 20)),
		std_logic_vector(to_signed(-829, 12) & to_signed(-449279, 20)),
		std_logic_vector(to_signed(-825, 12) & to_signed(-450106, 20)),
		std_logic_vector(to_signed(-821, 12) & to_signed(-450929, 20)),
		std_logic_vector(to_signed(-816, 12) & to_signed(-451747, 20)),
		std_logic_vector(to_signed(-812, 12) & to_signed(-452562, 20)),
		std_logic_vector(to_signed(-808, 12) & to_signed(-453372, 20)),
		std_logic_vector(to_signed(-804, 12) & to_signed(-454177, 20)),
		std_logic_vector(to_signed(-799, 12) & to_signed(-454979, 20)),
		std_logic_vector(to_signed(-795, 12) & to_signed(-455776, 20)),
		std_logic_vector(to_signed(-791, 12) & to_signed(-456569, 20)),
		std_logic_vector(to_signed(-786, 12) & to_signed(-457357, 20)),
		std_logic_vector(to_signed(-782, 12) & to_signed(-458141, 20)),
		std_logic_vector(to_signed(-778, 12) & to_signed(-458921, 20)),
		std_logic_vector(to_signed(-773, 12) & to_signed(-459697, 20)),
		std_logic_vector(to_signed(-769, 12) & to_signed(-460468, 20)),
		std_logic_vector(to_signed(-765, 12) & to_signed(-461235, 20)),
		std_logic_vector(to_signed(-760, 12) & to_signed(-461998, 20)),
		std_logic_vector(to_signed(-756, 12) & to_signed(-462756, 20)),
		std_logic_vector(to_signed(-752, 12) & to_signed(-463510, 20)),
		std_logic_vector(to_signed(-747, 12) & to_signed(-464259, 20)),
		std_logic_vector(to_signed(-743, 12) & to_signed(-465004, 20)),
		std_logic_vector(to_signed(-739, 12) & to_signed(-465745, 20)),
		std_logic_vector(to_signed(-734, 12) & to_signed(-466481, 20)),
		std_logic_vector(to_signed(-730, 12) & to_signed(-467213, 20)),
		std_logic_vector(to_signed(-725, 12) & to_signed(-467941, 20)),
		std_logic_vector(to_signed(-721, 12) & to_signed(-468664, 20)),
		std_logic_vector(to_signed(-717, 12) & to_signed(-469383, 20)),
		std_logic_vector(to_signed(-712, 12) & to_signed(-470097, 20)),
		std_logic_vector(to_signed(-708, 12) & to_signed(-470807, 20)),
		std_logic_vector(to_signed(-703, 12) & to_signed(-471513, 20)),
		std_logic_vector(to_signed(-699, 12) & to_signed(-472214, 20)),
		std_logic_vector(to_signed(-694, 12) & to_signed(-472911, 20)),
		std_logic_vector(to_signed(-690, 12) & to_signed(-473603, 20)),
		std_logic_vector(to_signed(-685, 12) & to_signed(-474290, 20)),
		std_logic_vector(to_signed(-681, 12) & to_signed(-474974, 20)),
		std_logic_vector(to_signed(-677, 12) & to_signed(-475652, 20)),
		std_logic_vector(to_signed(-672, 12) & to_signed(-476327, 20)),
		std_logic_vector(to_signed(-668, 12) & to_signed(-476997, 20)),
		std_logic_vector(to_signed(-663, 12) & to_signed(-477662, 20)),
		std_logic_vector(to_signed(-659, 12) & to_signed(-478323, 20)),
		std_logic_vector(to_signed(-654, 12) & to_signed(-478979, 20)),
		std_logic_vector(to_signed(-650, 12) & to_signed(-479631, 20)),
		std_logic_vector(to_signed(-645, 12) & to_signed(-480278, 20)),
		std_logic_vector(to_signed(-641, 12) & to_signed(-480921, 20)),
		std_logic_vector(to_signed(-636, 12) & to_signed(-481559, 20)),
		std_logic_vector(to_signed(-631, 12) & to_signed(-482193, 20)),
		std_logic_vector(to_signed(-627, 12) & to_signed(-482822, 20)),
		std_logic_vector(to_signed(-622, 12) & to_signed(-483447, 20)),
		std_logic_vector(to_signed(-618, 12) & to_signed(-484067, 20)),
		std_logic_vector(to_signed(-613, 12) & to_signed(-484682, 20)),
		std_logic_vector(to_signed(-609, 12) & to_signed(-485293, 20)),
		std_logic_vector(to_signed(-604, 12) & to_signed(-485900, 20)),
		std_logic_vector(to_signed(-600, 12) & to_signed(-486502, 20)),
		std_logic_vector(to_signed(-595, 12) & to_signed(-487099, 20)),
		std_logic_vector(to_signed(-590, 12) & to_signed(-487692, 20)),
		std_logic_vector(to_signed(-586, 12) & to_signed(-488280, 20)),
		std_logic_vector(to_signed(-581, 12) & to_signed(-488863, 20)),
		std_logic_vector(to_signed(-577, 12) & to_signed(-489442, 20)),
		std_logic_vector(to_signed(-572, 12) & to_signed(-490016, 20)),
		std_logic_vector(to_signed(-567, 12) & to_signed(-490586, 20)),
		std_logic_vector(to_signed(-563, 12) & to_signed(-491151, 20)),
		std_logic_vector(to_signed(-558, 12) & to_signed(-491711, 20)),
		std_logic_vector(to_signed(-553, 12) & to_signed(-492267, 20)),
		std_logic_vector(to_signed(-549, 12) & to_signed(-492818, 20)),
		std_logic_vector(to_signed(-544, 12) & to_signed(-493365, 20)),
		std_logic_vector(to_signed(-540, 12) & to_signed(-493907, 20)),
		std_logic_vector(to_signed(-535, 12) & to_signed(-494444, 20)),
		std_logic_vector(to_signed(-530, 12) & to_signed(-494977, 20)),
		std_logic_vector(to_signed(-526, 12) & to_signed(-495505, 20)),
		std_logic_vector(to_signed(-521, 12) & to_signed(-496028, 20)),
		std_logic_vector(to_signed(-516, 12) & to_signed(-496546, 20)),
		std_logic_vector(to_signed(-512, 12) & to_signed(-497060, 20)),
		std_logic_vector(to_signed(-507, 12) & to_signed(-497570, 20)),
		std_logic_vector(to_signed(-502, 12) & to_signed(-498074, 20)),
		std_logic_vector(to_signed(-498, 12) & to_signed(-498574, 20)),
		std_logic_vector(to_signed(-493, 12) & to_signed(-499069, 20)),
		std_logic_vector(to_signed(-488, 12) & to_signed(-499560, 20)),
		std_logic_vector(to_signed(-483, 12) & to_signed(-500045, 20)),
		std_logic_vector(to_signed(-479, 12) & to_signed(-500526, 20)),
		std_logic_vector(to_signed(-474, 12) & to_signed(-501003, 20)),
		std_logic_vector(to_signed(-469, 12) & to_signed(-501474, 20)),
		std_logic_vector(to_signed(-465, 12) & to_signed(-501941, 20)),
		std_logic_vector(to_signed(-460, 12) & to_signed(-502404, 20)),
		std_logic_vector(to_signed(-455, 12) & to_signed(-502861, 20)),
		std_logic_vector(to_signed(-450, 12) & to_signed(-503314, 20)),
		std_logic_vector(to_signed(-446, 12) & to_signed(-503762, 20)),
		std_logic_vector(to_signed(-441, 12) & to_signed(-504205, 20)),
		std_logic_vector(to_signed(-436, 12) & to_signed(-504644, 20)),
		std_logic_vector(to_signed(-431, 12) & to_signed(-505077, 20)),
		std_logic_vector(to_signed(-427, 12) & to_signed(-505506, 20)),
		std_logic_vector(to_signed(-422, 12) & to_signed(-505931, 20)),
		std_logic_vector(to_signed(-417, 12) & to_signed(-506350, 20)),
		std_logic_vector(to_signed(-412, 12) & to_signed(-506765, 20)),
		std_logic_vector(to_signed(-408, 12) & to_signed(-507175, 20)),
		std_logic_vector(to_signed(-403, 12) & to_signed(-507580, 20)),
		std_logic_vector(to_signed(-398, 12) & to_signed(-507980, 20)),
		std_logic_vector(to_signed(-393, 12) & to_signed(-508376, 20)),
		std_logic_vector(to_signed(-388, 12) & to_signed(-508767, 20)),
		std_logic_vector(to_signed(-384, 12) & to_signed(-509153, 20)),
		std_logic_vector(to_signed(-379, 12) & to_signed(-509534, 20)),
		std_logic_vector(to_signed(-374, 12) & to_signed(-509910, 20)),
		std_logic_vector(to_signed(-369, 12) & to_signed(-510282, 20)),
		std_logic_vector(to_signed(-364, 12) & to_signed(-510649, 20)),
		std_logic_vector(to_signed(-360, 12) & to_signed(-511011, 20)),
		std_logic_vector(to_signed(-355, 12) & to_signed(-511368, 20)),
		std_logic_vector(to_signed(-350, 12) & to_signed(-511721, 20)),
		std_logic_vector(to_signed(-345, 12) & to_signed(-512068, 20)),
		std_logic_vector(to_signed(-340, 12) & to_signed(-512411, 20)),
		std_logic_vector(to_signed(-336, 12) & to_signed(-512749, 20)),
		std_logic_vector(to_signed(-331, 12) & to_signed(-513082, 20)),
		std_logic_vector(to_signed(-326, 12) & to_signed(-513410, 20)),
		std_logic_vector(to_signed(-321, 12) & to_signed(-513734, 20)),
		std_logic_vector(to_signed(-316, 12) & to_signed(-514053, 20)),
		std_logic_vector(to_signed(-311, 12) & to_signed(-514366, 20)),
		std_logic_vector(to_signed(-307, 12) & to_signed(-514675, 20)),
		std_logic_vector(to_signed(-302, 12) & to_signed(-514979, 20)),
		std_logic_vector(to_signed(-297, 12) & to_signed(-515279, 20)),
		std_logic_vector(to_signed(-292, 12) & to_signed(-515573, 20)),
		std_logic_vector(to_signed(-287, 12) & to_signed(-515863, 20)),
		std_logic_vector(to_signed(-282, 12) & to_signed(-516147, 20)),
		std_logic_vector(to_signed(-277, 12) & to_signed(-516427, 20)),
		std_logic_vector(to_signed(-273, 12) & to_signed(-516702, 20)),
		std_logic_vector(to_signed(-268, 12) & to_signed(-516972, 20)),
		std_logic_vector(to_signed(-263, 12) & to_signed(-517238, 20)),
		std_logic_vector(to_signed(-258, 12) & to_signed(-517498, 20)),
		std_logic_vector(to_signed(-253, 12) & to_signed(-517753, 20)),
		std_logic_vector(to_signed(-248, 12) & to_signed(-518004, 20)),
		std_logic_vector(to_signed(-243, 12) & to_signed(-518250, 20)),
		std_logic_vector(to_signed(-238, 12) & to_signed(-518491, 20)),
		std_logic_vector(to_signed(-234, 12) & to_signed(-518727, 20)),
		std_logic_vector(to_signed(-229, 12) & to_signed(-518958, 20)),
		std_logic_vector(to_signed(-224, 12) & to_signed(-519184, 20)),
		std_logic_vector(to_signed(-219, 12) & to_signed(-519406, 20)),
		std_logic_vector(to_signed(-214, 12) & to_signed(-519622, 20)),
		std_logic_vector(to_signed(-209, 12) & to_signed(-519834, 20)),
		std_logic_vector(to_signed(-204, 12) & to_signed(-520040, 20)),
		std_logic_vector(to_signed(-199, 12) & to_signed(-520242, 20)),
		std_logic_vector(to_signed(-194, 12) & to_signed(-520439, 20)),
		std_logic_vector(to_signed(-190, 12) & to_signed(-520631, 20)),
		std_logic_vector(to_signed(-185, 12) & to_signed(-520818, 20)),
		std_logic_vector(to_signed(-180, 12) & to_signed(-521000, 20)),
		std_logic_vector(to_signed(-175, 12) & to_signed(-521178, 20)),
		std_logic_vector(to_signed(-170, 12) & to_signed(-521350, 20)),
		std_logic_vector(to_signed(-165, 12) & to_signed(-521517, 20)),
		std_logic_vector(to_signed(-160, 12) & to_signed(-521680, 20)),
		std_logic_vector(to_signed(-155, 12) & to_signed(-521838, 20)),
		std_logic_vector(to_signed(-150, 12) & to_signed(-521990, 20)),
		std_logic_vector(to_signed(-145, 12) & to_signed(-522138, 20)),
		std_logic_vector(to_signed(-140, 12) & to_signed(-522281, 20)),
		std_logic_vector(to_signed(-136, 12) & to_signed(-522419, 20)),
		std_logic_vector(to_signed(-131, 12) & to_signed(-522552, 20)),
		std_logic_vector(to_signed(-126, 12) & to_signed(-522680, 20)),
		std_logic_vector(to_signed(-121, 12) & to_signed(-522804, 20)),
		std_logic_vector(to_signed(-116, 12) & to_signed(-522922, 20)),
		std_logic_vector(to_signed(-111, 12) & to_signed(-523035, 20)),
		std_logic_vector(to_signed(-106, 12) & to_signed(-523144, 20)),
		std_logic_vector(to_signed(-101, 12) & to_signed(-523247, 20)),
		std_logic_vector(to_signed(-96, 12) & to_signed(-523346, 20)),
		std_logic_vector(to_signed(-91, 12) & to_signed(-523440, 20)),
		std_logic_vector(to_signed(-86, 12) & to_signed(-523529, 20)),
		std_logic_vector(to_signed(-81, 12) & to_signed(-523612, 20)),
		std_logic_vector(to_signed(-76, 12) & to_signed(-523691, 20)),
		std_logic_vector(to_signed(-72, 12) & to_signed(-523765, 20)),
		std_logic_vector(to_signed(-67, 12) & to_signed(-523834, 20)),
		std_logic_vector(to_signed(-62, 12) & to_signed(-523899, 20)),
		std_logic_vector(to_signed(-57, 12) & to_signed(-523958, 20)),
		std_logic_vector(to_signed(-52, 12) & to_signed(-524012, 20)),
		std_logic_vector(to_signed(-47, 12) & to_signed(-524061, 20)),
		std_logic_vector(to_signed(-42, 12) & to_signed(-524106, 20)),
		std_logic_vector(to_signed(-37, 12) & to_signed(-524145, 20)),
		std_logic_vector(to_signed(-32, 12) & to_signed(-524180, 20)),
		std_logic_vector(to_signed(-27, 12) & to_signed(-524209, 20)),
		std_logic_vector(to_signed(-22, 12) & to_signed(-524234, 20)),
		std_logic_vector(to_signed(-17, 12) & to_signed(-524254, 20)),
		std_logic_vector(to_signed(-12, 12) & to_signed(-524269, 20)),
		std_logic_vector(to_signed(-7, 12) & to_signed(-524278, 20)),
		std_logic_vector(to_signed(-2, 12) & to_signed(-524283, 20)),
		std_logic_vector(to_signed(2, 12) & to_signed(-524283, 20)),
		std_logic_vector(to_signed(7, 12) & to_signed(-524278, 20)),
		std_logic_vector(to_signed(12, 12) & to_signed(-524269, 20)),
		std_logic_vector(to_signed(17, 12) & to_signed(-524254, 20)),
		std_logic_vector(to_signed(22, 12) & to_signed(-524234, 20)),
		std_logic_vector(to_signed(27, 12) & to_signed(-524209, 20)),
		std_logic_vector(to_signed(32, 12) & to_signed(-524180, 20)),
		std_logic_vector(to_signed(37, 12) & to_signed(-524145, 20)),
		std_logic_vector(to_signed(42, 12) & to_signed(-524106, 20)),
		std_logic_vector(to_signed(47, 12) & to_signed(-524061, 20)),
		std_logic_vector(to_signed(52, 12) & to_signed(-524012, 20)),
		std_logic_vector(to_signed(57, 12) & to_signed(-523958, 20)),
		std_logic_vector(to_signed(62, 12) & to_signed(-523899, 20)),
		std_logic_vector(to_signed(67, 12) & to_signed(-523834, 20)),
		std_logic_vector(to_signed(72, 12) & to_signed(-523765, 20)),
		std_logic_vector(to_signed(76, 12) & to_signed(-523691, 20)),
		std_logic_vector(to_signed(81, 12) & to_signed(-523612, 20)),
		std_logic_vector(to_signed(86, 12) & to_signed(-523529, 20)),
		std_logic_vector(to_signed(91, 12) & to_signed(-523440, 20)),
		std_logic_vector(to_signed(96, 12) & to_signed(-523346, 20)),
		std_logic_vector(to_signed(101, 12) & to_signed(-523247, 20)),
		std_logic_vector(to_signed(106, 12) & to_signed(-523144, 20)),
		std_logic_vector(to_signed(111, 12) & to_signed(-523035, 20)),
		std_logic_vector(to_signed(116, 12) & to_signed(-522922, 20)),
		std_logic_vector(to_signed(121, 12) & to_signed(-522804, 20)),
		std_logic_vector(to_signed(126, 12) & to_signed(-522680, 20)),
		std_logic_vector(to_signed(131, 12) & to_signed(-522552, 20)),
		std_logic_vector(to_signed(136, 12) & to_signed(-522419, 20)),
		std_logic_vector(to_signed(140, 12) & to_signed(-522281, 20)),
		std_logic_vector(to_signed(145, 12) & to_signed(-522138, 20)),
		std_logic_vector(to_signed(150, 12) & to_signed(-521990, 20)),
		std_logic_vector(to_signed(155, 12) & to_signed(-521838, 20)),
		std_logic_vector(to_signed(160, 12) & to_signed(-521680, 20)),
		std_logic_vector(to_signed(165, 12) & to_signed(-521517, 20)),
		std_logic_vector(to_signed(170, 12) & to_signed(-521350, 20)),
		std_logic_vector(to_signed(175, 12) & to_signed(-521178, 20)),
		std_logic_vector(to_signed(180, 12) & to_signed(-521000, 20)),
		std_logic_vector(to_signed(185, 12) & to_signed(-520818, 20)),
		std_logic_vector(to_signed(190, 12) & to_signed(-520631, 20)),
		std_logic_vector(to_signed(194, 12) & to_signed(-520439, 20)),
		std_logic_vector(to_signed(199, 12) & to_signed(-520242, 20)),
		std_logic_vector(to_signed(204, 12) & to_signed(-520040, 20)),
		std_logic_vector(to_signed(209, 12) & to_signed(-519834, 20)),
		std_logic_vector(to_signed(214, 12) & to_signed(-519622, 20)),
		std_logic_vector(to_signed(219, 12) & to_signed(-519406, 20)),
		std_logic_vector(to_signed(224, 12) & to_signed(-519184, 20)),
		std_logic_vector(to_signed(229, 12) & to_signed(-518958, 20)),
		std_logic_vector(to_signed(234, 12) & to_signed(-518727, 20)),
		std_logic_vector(to_signed(238, 12) & to_signed(-518491, 20)),
		std_logic_vector(to_signed(243, 12) & to_signed(-518250, 20)),
		std_logic_vector(to_signed(248, 12) & to_signed(-518004, 20)),
		std_logic_vector(to_signed(253, 12) & to_signed(-517753, 20)),
		std_logic_vector(to_signed(258, 12) & to_signed(-517498, 20)),
		std_logic_vector(to_signed(263, 12) & to_signed(-517238, 20)),
		std_logic_vector(to_signed(268, 12) & to_signed(-516972, 20)),
		std_logic_vector(to_signed(273, 12) & to_signed(-516702, 20)),
		std_logic_vector(to_signed(277, 12) & to_signed(-516427, 20)),
		std_logic_vector(to_signed(282, 12) & to_signed(-516147, 20)),
		std_logic_vector(to_signed(287, 12) & to_signed(-515863, 20)),
		std_logic_vector(to_signed(292, 12) & to_signed(-515573, 20)),
		std_logic_vector(to_signed(297, 12) & to_signed(-515279, 20)),
		std_logic_vector(to_signed(302, 12) & to_signed(-514979, 20)),
		std_logic_vector(to_signed(307, 12) & to_signed(-514675, 20)),
		std_logic_vector(to_signed(311, 12) & to_signed(-514366, 20)),
		std_logic_vector(to_signed(316, 12) & to_signed(-514053, 20)),
		std_logic_vector(to_signed(321, 12) & to_signed(-513734, 20)),
		std_logic_vector(to_signed(326, 12) & to_signed(-513410, 20)),
		std_logic_vector(to_signed(331, 12) & to_signed(-513082, 20)),
		std_logic_vector(to_signed(336, 12) & to_signed(-512749, 20)),
		std_logic_vector(to_signed(340, 12) & to_signed(-512411, 20)),
		std_logic_vector(to_signed(345, 12) & to_signed(-512068, 20)),
		std_logic_vector(to_signed(350, 12) & to_signed(-511721, 20)),
		std_logic_vector(to_signed(355, 12) & to_signed(-511368, 20)),
		std_logic_vector(to_signed(360, 12) & to_signed(-511011, 20)),
		std_logic_vector(to_signed(364, 12) & to_signed(-510649, 20)),
		std_logic_vector(to_signed(369, 12) & to_signed(-510282, 20)),
		std_logic_vector(to_signed(374, 12) & to_signed(-509910, 20)),
		std_logic_vector(to_signed(379, 12) & to_signed(-509534, 20)),
		std_logic_vector(to_signed(384, 12) & to_signed(-509153, 20)),
		std_logic_vector(to_signed(388, 12) & to_signed(-508767, 20)),
		std_logic_vector(to_signed(393, 12) & to_signed(-508376, 20)),
		std_logic_vector(to_signed(398, 12) & to_signed(-507980, 20)),
		std_logic_vector(to_signed(403, 12) & to_signed(-507580, 20)),
		std_logic_vector(to_signed(408, 12) & to_signed(-507175, 20)),
		std_logic_vector(to_signed(412, 12) & to_signed(-506765, 20)),
		std_logic_vector(to_signed(417, 12) & to_signed(-506350, 20)),
		std_logic_vector(to_signed(422, 12) & to_signed(-505931, 20)),
		std_logic_vector(to_signed(427, 12) & to_signed(-505506, 20)),
		std_logic_vector(to_signed(431, 12) & to_signed(-505077, 20)),
		std_logic_vector(to_signed(436, 12) & to_signed(-504644, 20)),
		std_logic_vector(to_signed(441, 12) & to_signed(-504205, 20)),
		std_logic_vector(to_signed(446, 12) & to_signed(-503762, 20)),
		std_logic_vector(to_signed(450, 12) & to_signed(-503314, 20)),
		std_logic_vector(to_signed(455, 12) & to_signed(-502861, 20)),
		std_logic_vector(to_signed(460, 12) & to_signed(-502404, 20)),
		std_logic_vector(to_signed(465, 12) & to_signed(-501941, 20)),
		std_logic_vector(to_signed(469, 12) & to_signed(-501474, 20)),
		std_logic_vector(to_signed(474, 12) & to_signed(-501003, 20)),
		std_logic_vector(to_signed(479, 12) & to_signed(-500526, 20)),
		std_logic_vector(to_signed(483, 12) & to_signed(-500045, 20)),
		std_logic_vector(to_signed(488, 12) & to_signed(-499560, 20)),
		std_logic_vector(to_signed(493, 12) & to_signed(-499069, 20)),
		std_logic_vector(to_signed(498, 12) & to_signed(-498574, 20)),
		std_logic_vector(to_signed(502, 12) & to_signed(-498074, 20)),
		std_logic_vector(to_signed(507, 12) & to_signed(-497570, 20)),
		std_logic_vector(to_signed(512, 12) & to_signed(-497060, 20)),
		std_logic_vector(to_signed(516, 12) & to_signed(-496546, 20)),
		std_logic_vector(to_signed(521, 12) & to_signed(-496028, 20)),
		std_logic_vector(to_signed(526, 12) & to_signed(-495505, 20)),
		std_logic_vector(to_signed(530, 12) & to_signed(-494977, 20)),
		std_logic_vector(to_signed(535, 12) & to_signed(-494444, 20)),
		std_logic_vector(to_signed(540, 12) & to_signed(-493907, 20)),
		std_logic_vector(to_signed(544, 12) & to_signed(-493365, 20)),
		std_logic_vector(to_signed(549, 12) & to_signed(-492818, 20)),
		std_logic_vector(to_signed(553, 12) & to_signed(-492267, 20)),
		std_logic_vector(to_signed(558, 12) & to_signed(-491711, 20)),
		std_logic_vector(to_signed(563, 12) & to_signed(-491151, 20)),
		std_logic_vector(to_signed(567, 12) & to_signed(-490586, 20)),
		std_logic_vector(to_signed(572, 12) & to_signed(-490016, 20)),
		std_logic_vector(to_signed(577, 12) & to_signed(-489442, 20)),
		std_logic_vector(to_signed(581, 12) & to_signed(-488863, 20)),
		std_logic_vector(to_signed(586, 12) & to_signed(-488280, 20)),
		std_logic_vector(to_signed(590, 12) & to_signed(-487692, 20)),
		std_logic_vector(to_signed(595, 12) & to_signed(-487099, 20)),
		std_logic_vector(to_signed(600, 12) & to_signed(-486502, 20)),
		std_logic_vector(to_signed(604, 12) & to_signed(-485900, 20)),
		std_logic_vector(to_signed(609, 12) & to_signed(-485293, 20)),
		std_logic_vector(to_signed(613, 12) & to_signed(-484682, 20)),
		std_logic_vector(to_signed(618, 12) & to_signed(-484067, 20)),
		std_logic_vector(to_signed(622, 12) & to_signed(-483447, 20)),
		std_logic_vector(to_signed(627, 12) & to_signed(-482822, 20)),
		std_logic_vector(to_signed(631, 12) & to_signed(-482193, 20)),
		std_logic_vector(to_signed(636, 12) & to_signed(-481559, 20)),
		std_logic_vector(to_signed(641, 12) & to_signed(-480921, 20)),
		std_logic_vector(to_signed(645, 12) & to_signed(-480278, 20)),
		std_logic_vector(to_signed(650, 12) & to_signed(-479631, 20)),
		std_logic_vector(to_signed(654, 12) & to_signed(-478979, 20)),
		std_logic_vector(to_signed(659, 12) & to_signed(-478323, 20)),
		std_logic_vector(to_signed(663, 12) & to_signed(-477662, 20)),
		std_logic_vector(to_signed(668, 12) & to_signed(-476997, 20)),
		std_logic_vector(to_signed(672, 12) & to_signed(-476327, 20)),
		std_logic_vector(to_signed(677, 12) & to_signed(-475652, 20)),
		std_logic_vector(to_signed(681, 12) & to_signed(-474974, 20)),
		std_logic_vector(to_signed(685, 12) & to_signed(-474290, 20)),
		std_logic_vector(to_signed(690, 12) & to_signed(-473603, 20)),
		std_logic_vector(to_signed(694, 12) & to_signed(-472911, 20)),
		std_logic_vector(to_signed(699, 12) & to_signed(-472214, 20)),
		std_logic_vector(to_signed(703, 12) & to_signed(-471513, 20)),
		std_logic_vector(to_signed(708, 12) & to_signed(-470807, 20)),
		std_logic_vector(to_signed(712, 12) & to_signed(-470097, 20)),
		std_logic_vector(to_signed(717, 12) & to_signed(-469383, 20)),
		std_logic_vector(to_signed(721, 12) & to_signed(-468664, 20)),
		std_logic_vector(to_signed(725, 12) & to_signed(-467941, 20)),
		std_logic_vector(to_signed(730, 12) & to_signed(-467213, 20)),
		std_logic_vector(to_signed(734, 12) & to_signed(-466481, 20)),
		std_logic_vector(to_signed(739, 12) & to_signed(-465745, 20)),
		std_logic_vector(to_signed(743, 12) & to_signed(-465004, 20)),
		std_logic_vector(to_signed(747, 12) & to_signed(-464259, 20)),
		std_logic_vector(to_signed(752, 12) & to_signed(-463510, 20)),
		std_logic_vector(to_signed(756, 12) & to_signed(-462756, 20)),
		std_logic_vector(to_signed(760, 12) & to_signed(-461998, 20)),
		std_logic_vector(to_signed(765, 12) & to_signed(-461235, 20)),
		std_logic_vector(to_signed(769, 12) & to_signed(-460468, 20)),
		std_logic_vector(to_signed(773, 12) & to_signed(-459697, 20)),
		std_logic_vector(to_signed(778, 12) & to_signed(-458921, 20)),
		std_logic_vector(to_signed(782, 12) & to_signed(-458141, 20)),
		std_logic_vector(to_signed(786, 12) & to_signed(-457357, 20)),
		std_logic_vector(to_signed(791, 12) & to_signed(-456569, 20)),
		std_logic_vector(to_signed(795, 12) & to_signed(-455776, 20)),
		std_logic_vector(to_signed(799, 12) & to_signed(-454979, 20)),
		std_logic_vector(to_signed(804, 12) & to_signed(-454177, 20)),
		std_logic_vector(to_signed(808, 12) & to_signed(-453372, 20)),
		std_logic_vector(to_signed(812, 12) & to_signed(-452562, 20)),
		std_logic_vector(to_signed(816, 12) & to_signed(-451747, 20)),
		std_logic_vector(to_signed(821, 12) & to_signed(-450929, 20)),
		std_logic_vector(to_signed(825, 12) & to_signed(-450106, 20)),
		std_logic_vector(to_signed(829, 12) & to_signed(-449279, 20)),
		std_logic_vector(to_signed(833, 12) & to_signed(-448448, 20)),
		std_logic_vector(to_signed(837, 12) & to_signed(-447613, 20)),
		std_logic_vector(to_signed(842, 12) & to_signed(-446773, 20)),
		std_logic_vector(to_signed(846, 12) & to_signed(-445929, 20)),
		std_logic_vector(to_signed(850, 12) & to_signed(-445081, 20)),
		std_logic_vector(to_signed(854, 12) & to_signed(-444229, 20)),
		std_logic_vector(to_signed(858, 12) & to_signed(-443373, 20)),
		std_logic_vector(to_signed(863, 12) & to_signed(-442512, 20)),
		std_logic_vector(to_signed(867, 12) & to_signed(-441648, 20)),
		std_logic_vector(to_signed(871, 12) & to_signed(-440779, 20)),
		std_logic_vector(to_signed(875, 12) & to_signed(-439906, 20)),
		std_logic_vector(to_signed(879, 12) & to_signed(-439029, 20)),
		std_logic_vector(to_signed(883, 12) & to_signed(-438147, 20)),
		std_logic_vector(to_signed(887, 12) & to_signed(-437262, 20)),
		std_logic_vector(to_signed(892, 12) & to_signed(-436373, 20)),
		std_logic_vector(to_signed(896, 12) & to_signed(-435479, 20)),
		std_logic_vector(to_signed(900, 12) & to_signed(-434581, 20)),
		std_logic_vector(to_signed(904, 12) & to_signed(-433679, 20)),
		std_logic_vector(to_signed(908, 12) & to_signed(-432773, 20)),
		std_logic_vector(to_signed(912, 12) & to_signed(-431863, 20)),
		std_logic_vector(to_signed(916, 12) & to_signed(-430949, 20)),
		std_logic_vector(to_signed(920, 12) & to_signed(-430031, 20)),
		std_logic_vector(to_signed(924, 12) & to_signed(-429109, 20)),
		std_logic_vector(to_signed(928, 12) & to_signed(-428183, 20)),
		std_logic_vector(to_signed(932, 12) & to_signed(-427253, 20)),
		std_logic_vector(to_signed(936, 12) & to_signed(-426319, 20)),
		std_logic_vector(to_signed(940, 12) & to_signed(-425380, 20)),
		std_logic_vector(to_signed(944, 12) & to_signed(-424438, 20)),
		std_logic_vector(to_signed(948, 12) & to_signed(-423492, 20)),
		std_logic_vector(to_signed(952, 12) & to_signed(-422542, 20)),
		std_logic_vector(to_signed(956, 12) & to_signed(-421587, 20)),
		std_logic_vector(to_signed(960, 12) & to_signed(-420629, 20)),
		std_logic_vector(to_signed(964, 12) & to_signed(-419667, 20)),
		std_logic_vector(to_signed(968, 12) & to_signed(-418701, 20)),
		std_logic_vector(to_signed(972, 12) & to_signed(-417731, 20)),
		std_logic_vector(to_signed(976, 12) & to_signed(-416757, 20)),
		std_logic_vector(to_signed(980, 12) & to_signed(-415779, 20)),
		std_logic_vector(to_signed(984, 12) & to_signed(-414797, 20)),
		std_logic_vector(to_signed(988, 12) & to_signed(-413812, 20)),
		std_logic_vector(to_signed(992, 12) & to_signed(-412822, 20)),
		std_logic_vector(to_signed(995, 12) & to_signed(-411829, 20)),
		std_logic_vector(to_signed(999, 12) & to_signed(-410831, 20)),
		std_logic_vector(to_signed(1003, 12) & to_signed(-409830, 20)),
		std_logic_vector(to_signed(1007, 12) & to_signed(-408825, 20)),
		std_logic_vector(to_signed(1011, 12) & to_signed(-407816, 20)),
		std_logic_vector(to_signed(1015, 12) & to_signed(-406803, 20)),
		std_logic_vector(to_signed(1019, 12) & to_signed(-405787, 20)),
		std_logic_vector(to_signed(1022, 12) & to_signed(-404766, 20)),
		std_logic_vector(to_signed(1026, 12) & to_signed(-403742, 20)),
		std_logic_vector(to_signed(1030, 12) & to_signed(-402714, 20)),
		std_logic_vector(to_signed(1034, 12) & to_signed(-401682, 20)),
		std_logic_vector(to_signed(1037, 12) & to_signed(-400647, 20)),
		std_logic_vector(to_signed(1041, 12) & to_signed(-399607, 20)),
		std_logic_vector(to_signed(1045, 12) & to_signed(-398564, 20)),
		std_logic_vector(to_signed(1049, 12) & to_signed(-397517, 20)),
		std_logic_vector(to_signed(1052, 12) & to_signed(-396467, 20)),
		std_logic_vector(to_signed(1056, 12) & to_signed(-395412, 20)),
		std_logic_vector(to_signed(1060, 12) & to_signed(-394354, 20)),
		std_logic_vector(to_signed(1064, 12) & to_signed(-393293, 20)),
		std_logic_vector(to_signed(1067, 12) & to_signed(-392227, 20)),
		std_logic_vector(to_signed(1071, 12) & to_signed(-391158, 20)),
		std_logic_vector(to_signed(1075, 12) & to_signed(-390085, 20)),
		std_logic_vector(to_signed(1078, 12) & to_signed(-389008, 20)),
		std_logic_vector(to_signed(1082, 12) & to_signed(-387928, 20)),
		std_logic_vector(to_signed(1086, 12) & to_signed(-386844, 20)),
		std_logic_vector(to_signed(1089, 12) & to_signed(-385757, 20)),
		std_logic_vector(to_signed(1093, 12) & to_signed(-384666, 20)),
		std_logic_vector(to_signed(1097, 12) & to_signed(-383571, 20)),
		std_logic_vector(to_signed(1100, 12) & to_signed(-382473, 20)),
		std_logic_vector(to_signed(1104, 12) & to_signed(-381371, 20)),
		std_logic_vector(to_signed(1107, 12) & to_signed(-380265, 20)),
		std_logic_vector(to_signed(1111, 12) & to_signed(-379156, 20)),
		std_logic_vector(to_signed(1114, 12) & to_signed(-378043, 20)),
		std_logic_vector(to_signed(1118, 12) & to_signed(-376927, 20)),
		std_logic_vector(to_signed(1122, 12) & to_signed(-375807, 20)),
		std_logic_vector(to_signed(1125, 12) & to_signed(-374684, 20)),
		std_logic_vector(to_signed(1129, 12) & to_signed(-373557, 20)),
		std_logic_vector(to_signed(1132, 12) & to_signed(-372427, 20)),
		std_logic_vector(to_signed(1136, 12) & to_signed(-371293, 20)),
		std_logic_vector(to_signed(1139, 12) & to_signed(-370156, 20)),
		std_logic_vector(to_signed(1143, 12) & to_signed(-369015, 20)),
		std_logic_vector(to_signed(1146, 12) & to_signed(-367870, 20)),
		std_logic_vector(to_signed(1150, 12) & to_signed(-366723, 20)),
		std_logic_vector(to_signed(1153, 12) & to_signed(-365571, 20)),
		std_logic_vector(to_signed(1156, 12) & to_signed(-364417, 20)),
		std_logic_vector(to_signed(1160, 12) & to_signed(-363259, 20)),
		std_logic_vector(to_signed(1163, 12) & to_signed(-362097, 20)),
		std_logic_vector(to_signed(1167, 12) & to_signed(-360932, 20)),
		std_logic_vector(to_signed(1170, 12) & to_signed(-359764, 20)),
		std_logic_vector(to_signed(1173, 12) & to_signed(-358592, 20)),
		std_logic_vector(to_signed(1177, 12) & to_signed(-357417, 20)),
		std_logic_vector(to_signed(1180, 12) & to_signed(-356239, 20)),
		std_logic_vector(to_signed(1183, 12) & to_signed(-355057, 20)),
		std_logic_vector(to_signed(1187, 12) & to_signed(-353872, 20)),
		std_logic_vector(to_signed(1190, 12) & to_signed(-352683, 20)),
		std_logic_vector(to_signed(1193, 12) & to_signed(-351491, 20)),
		std_logic_vector(to_signed(1197, 12) & to_signed(-350296, 20)),
		std_logic_vector(to_signed(1200, 12) & to_signed(-349098, 20)),
		std_logic_vector(to_signed(1203, 12) & to_signed(-347896, 20)),
		std_logic_vector(to_signed(1207, 12) & to_signed(-346691, 20)),
		std_logic_vector(to_signed(1210, 12) & to_signed(-345483, 20)),
		std_logic_vector(to_signed(1213, 12) & to_signed(-344271, 20)),
		std_logic_vector(to_signed(1216, 12) & to_signed(-343057, 20)),
		std_logic_vector(to_signed(1220, 12) & to_signed(-341839, 20)),
		std_logic_vector(to_signed(1223, 12) & to_signed(-340618, 20)),
		std_logic_vector(to_signed(1226, 12) & to_signed(-339393, 20)),
		std_logic_vector(to_signed(1229, 12) & to_signed(-338166, 20)),
		std_logic_vector(to_signed(1232, 12) & to_signed(-336935, 20)),
		std_logic_vector(to_signed(1236, 12) & to_signed(-335701, 20)),
		std_logic_vector(to_signed(1239, 12) & to_signed(-334464, 20)),
		std_logic_vector(to_signed(1242, 12) & to_signed(-333224, 20)),
		std_logic_vector(to_signed(1245, 12) & to_signed(-331980, 20)),
		std_logic_vector(to_signed(1248, 12) & to_signed(-330734, 20)),
		std_logic_vector(to_signed(1251, 12) & to_signed(-329484, 20)),
		std_logic_vector(to_signed(1254, 12) & to_signed(-328231, 20)),
		std_logic_vector(to_signed(1257, 12) & to_signed(-326976, 20)),
		std_logic_vector(to_signed(1260, 12) & to_signed(-325717, 20)),
		std_logic_vector(to_signed(1263, 12) & to_signed(-324455, 20)),
		std_logic_vector(to_signed(1267, 12) & to_signed(-323190, 20)),
		std_logic_vector(to_signed(1270, 12) & to_signed(-321922, 20)),
		std_logic_vector(to_signed(1273, 12) & to_signed(-320651, 20)),
		std_logic_vector(to_signed(1276, 12) & to_signed(-319377, 20)),
		std_logic_vector(to_signed(1279, 12) & to_signed(-318099, 20)),
		std_logic_vector(to_signed(1282, 12) & to_signed(-316819, 20)),
		std_logic_vector(to_signed(1285, 12) & to_signed(-315536, 20)),
		std_logic_vector(to_signed(1288, 12) & to_signed(-314250, 20)),
		std_logic_vector(to_signed(1290, 12) & to_signed(-312961, 20)),
		std_logic_vector(to_signed(1293, 12) & to_signed(-311669, 20)),
		std_logic_vector(to_signed(1296, 12) & to_signed(-310374, 20)),
		std_logic_vector(to_signed(1299, 12) & to_signed(-309077, 20)),
		std_logic_vector(to_signed(1302, 12) & to_signed(-307776, 20)),
		std_logic_vector(to_signed(1305, 12) & to_signed(-306472, 20)),
		std_logic_vector(to_signed(1308, 12) & to_signed(-305166, 20)),
		std_logic_vector(to_signed(1311, 12) & to_signed(-303856, 20)),
		std_logic_vector(to_signed(1314, 12) & to_signed(-302544, 20)),
		std_logic_vector(to_signed(1316, 12) & to_signed(-301229, 20)),
		std_logic_vector(to_signed(1319, 12) & to_signed(-299911, 20)),
		std_logic_vector(to_signed(1322, 12) & to_signed(-298590, 20)),
		std_logic_vector(to_signed(1325, 12) & to_signed(-297267, 20)),
		std_logic_vector(to_signed(1328, 12) & to_signed(-295941, 20)),
		std_logic_vector(to_signed(1331, 12) & to_signed(-294611, 20)),
		std_logic_vector(to_signed(1333, 12) & to_signed(-293280, 20)),
		std_logic_vector(to_signed(1336, 12) & to_signed(-291945, 20)),
		std_logic_vector(to_signed(1339, 12) & to_signed(-290608, 20)),
		std_logic_vector(to_signed(1342, 12) & to_signed(-289267, 20)),
		std_logic_vector(to_signed(1344, 12) & to_signed(-287925, 20)),
		std_logic_vector(to_signed(1347, 12) & to_signed(-286579, 20)),
		std_logic_vector(to_signed(1350, 12) & to_signed(-285231, 20)),
		std_logic_vector(to_signed(1352, 12) & to_signed(-283880, 20)),
		std_logic_vector(to_signed(1355, 12) & to_signed(-282526, 20)),
		std_logic_vector(to_signed(1358, 12) & to_signed(-281170, 20)),
		std_logic_vector(to_signed(1360, 12) & to_signed(-279811, 20)),
		std_logic_vector(to_signed(1363, 12) & to_signed(-278449, 20)),
		std_logic_vector(to_signed(1365, 12) & to_signed(-277085, 20)),
		std_logic_vector(to_signed(1368, 12) & to_signed(-275718, 20)),
		std_logic_vector(to_signed(1371, 12) & to_signed(-274349, 20)),
		std_logic_vector(to_signed(1373, 12) & to_signed(-272977, 20)),
		std_logic_vector(to_signed(1376, 12) & to_signed(-271602, 20)),
		std_logic_vector(to_signed(1378, 12) & to_signed(-270225, 20)),
		std_logic_vector(to_signed(1381, 12) & to_signed(-268846, 20)),
		std_logic_vector(to_signed(1383, 12) & to_signed(-267464, 20)),
		std_logic_vector(to_signed(1386, 12) & to_signed(-266079, 20)),
		std_logic_vector(to_signed(1388, 12) & to_signed(-264692, 20)),
		std_logic_vector(to_signed(1391, 12) & to_signed(-263302, 20)),
		std_logic_vector(to_signed(1393, 12) & to_signed(-261910, 20)),
		std_logic_vector(to_signed(1396, 12) & to_signed(-260515, 20)),
		std_logic_vector(to_signed(1398, 12) & to_signed(-259118, 20)),
		std_logic_vector(to_signed(1401, 12) & to_signed(-257719, 20)),
		std_logic_vector(to_signed(1403, 12) & to_signed(-256317, 20)),
		std_logic_vector(to_signed(1406, 12) & to_signed(-254912, 20)),
		std_logic_vector(to_signed(1408, 12) & to_signed(-253506, 20)),
		std_logic_vector(to_signed(1410, 12) & to_signed(-252096, 20)),
		std_logic_vector(to_signed(1413, 12) & to_signed(-250685, 20)),
		std_logic_vector(to_signed(1415, 12) & to_signed(-249271, 20)),
		std_logic_vector(to_signed(1417, 12) & to_signed(-247855, 20)),
		std_logic_vector(to_signed(1420, 12) & to_signed(-246436, 20)),
		std_logic_vector(to_signed(1422, 12) & to_signed(-245015, 20)),
		std_logic_vector(to_signed(1424, 12) & to_signed(-243592, 20)),
		std_logic_vector(to_signed(1427, 12) & to_signed(-242167, 20)),
		std_logic_vector(to_signed(1429, 12) & to_signed(-240739, 20)),
		std_logic_vector(to_signed(1431, 12) & to_signed(-239309, 20)),
		std_logic_vector(to_signed(1433, 12) & to_signed(-237877, 20)),
		std_logic_vector(to_signed(1436, 12) & to_signed(-236442, 20)),
		std_logic_vector(to_signed(1438, 12) & to_signed(-235005, 20)),
		std_logic_vector(to_signed(1440, 12) & to_signed(-233566, 20)),
		std_logic_vector(to_signed(1442, 12) & to_signed(-232125, 20)),
		std_logic_vector(to_signed(1444, 12) & to_signed(-230682, 20)),
		std_logic_vector(to_signed(1447, 12) & to_signed(-229236, 20)),
		std_logic_vector(to_signed(1449, 12) & to_signed(-227789, 20)),
		std_logic_vector(to_signed(1451, 12) & to_signed(-226339, 20)),
		std_logic_vector(to_signed(1453, 12) & to_signed(-224887, 20)),
		std_logic_vector(to_signed(1455, 12) & to_signed(-223433, 20)),
		std_logic_vector(to_signed(1457, 12) & to_signed(-221977, 20)),
		std_logic_vector(to_signed(1459, 12) & to_signed(-220519, 20)),
		std_logic_vector(to_signed(1461, 12) & to_signed(-219058, 20)),
		std_logic_vector(to_signed(1463, 12) & to_signed(-217596, 20)),
		std_logic_vector(to_signed(1465, 12) & to_signed(-216131, 20)),
		std_logic_vector(to_signed(1467, 12) & to_signed(-214665, 20)),
		std_logic_vector(to_signed(1469, 12) & to_signed(-213197, 20)),
		std_logic_vector(to_signed(1471, 12) & to_signed(-211726, 20)),
		std_logic_vector(to_signed(1473, 12) & to_signed(-210254, 20)),
		std_logic_vector(to_signed(1475, 12) & to_signed(-208779, 20)),
		std_logic_vector(to_signed(1477, 12) & to_signed(-207303, 20)),
		std_logic_vector(to_signed(1479, 12) & to_signed(-205824, 20)),
		std_logic_vector(to_signed(1481, 12) & to_signed(-204344, 20)),
		std_logic_vector(to_signed(1483, 12) & to_signed(-202862, 20)),
		std_logic_vector(to_signed(1485, 12) & to_signed(-201378, 20)),
		std_logic_vector(to_signed(1487, 12) & to_signed(-199892, 20)),
		std_logic_vector(to_signed(1489, 12) & to_signed(-198404, 20)),
		std_logic_vector(to_signed(1491, 12) & to_signed(-196914, 20)),
		std_logic_vector(to_signed(1493, 12) & to_signed(-195422, 20)),
		std_logic_vector(to_signed(1494, 12) & to_signed(-193929, 20)),
		std_logic_vector(to_signed(1496, 12) & to_signed(-192433, 20)),
		std_logic_vector(to_signed(1498, 12) & to_signed(-190936, 20)),
		std_logic_vector(to_signed(1500, 12) & to_signed(-189437, 20)),
		std_logic_vector(to_signed(1502, 12) & to_signed(-187937, 20)),
		std_logic_vector(to_signed(1503, 12) & to_signed(-186434, 20)),
		std_logic_vector(to_signed(1505, 12) & to_signed(-184930, 20)),
		std_logic_vector(to_signed(1507, 12) & to_signed(-183424, 20)),
		std_logic_vector(to_signed(1509, 12) & to_signed(-181916, 20)),
		std_logic_vector(to_signed(1510, 12) & to_signed(-180407, 20)),
		std_logic_vector(to_signed(1512, 12) & to_signed(-178896, 20)),
		std_logic_vector(to_signed(1514, 12) & to_signed(-177383, 20)),
		std_logic_vector(to_signed(1515, 12) & to_signed(-175869, 20)),
		std_logic_vector(to_signed(1517, 12) & to_signed(-174352, 20)),
		std_logic_vector(to_signed(1519, 12) & to_signed(-172835, 20)),
		std_logic_vector(to_signed(1520, 12) & to_signed(-171315, 20)),
		std_logic_vector(to_signed(1522, 12) & to_signed(-169794, 20)),
		std_logic_vector(to_signed(1523, 12) & to_signed(-168272, 20)),
		std_logic_vector(to_signed(1525, 12) & to_signed(-166748, 20)),
		std_logic_vector(to_signed(1527, 12) & to_signed(-165222, 20)),
		std_logic_vector(to_signed(1528, 12) & to_signed(-163694, 20)),
		std_logic_vector(to_signed(1530, 12) & to_signed(-162166, 20)),
		std_logic_vector(to_signed(1531, 12) & to_signed(-160635, 20)),
		std_logic_vector(to_signed(1533, 12) & to_signed(-159103, 20)),
		std_logic_vector(to_signed(1534, 12) & to_signed(-157570, 20)),
		std_logic_vector(to_signed(1536, 12) & to_signed(-156035, 20)),
		std_logic_vector(to_signed(1537, 12) & to_signed(-154499, 20)),
		std_logic_vector(to_signed(1539, 12) & to_signed(-152961, 20)),
		std_logic_vector(to_signed(1540, 12) & to_signed(-151422, 20)),
		std_logic_vector(to_signed(1541, 12) & to_signed(-149881, 20)),
		std_logic_vector(to_signed(1543, 12) & to_signed(-148339, 20)),
		std_logic_vector(to_signed(1544, 12) & to_signed(-146796, 20)),
		std_logic_vector(to_signed(1546, 12) & to_signed(-145251, 20)),
		std_logic_vector(to_signed(1547, 12) & to_signed(-143705, 20)),
		std_logic_vector(to_signed(1548, 12) & to_signed(-142157, 20)),
		std_logic_vector(to_signed(1550, 12) & to_signed(-140608, 20)),
		std_logic_vector(to_signed(1551, 12) & to_signed(-139058, 20)),
		std_logic_vector(to_signed(1552, 12) & to_signed(-137506, 20)),
		std_logic_vector(to_signed(1553, 12) & to_signed(-135954, 20)),
		std_logic_vector(to_signed(1555, 12) & to_signed(-134400, 20)),
		std_logic_vector(to_signed(1556, 12) & to_signed(-132844, 20)),
		std_logic_vector(to_signed(1557, 12) & to_signed(-131288, 20)),
		std_logic_vector(to_signed(1558, 12) & to_signed(-129730, 20)),
		std_logic_vector(to_signed(1560, 12) & to_signed(-128171, 20)),
		std_logic_vector(to_signed(1561, 12) & to_signed(-126610, 20)),
		std_logic_vector(to_signed(1562, 12) & to_signed(-125049, 20)),
		std_logic_vector(to_signed(1563, 12) & to_signed(-123486, 20)),
		std_logic_vector(to_signed(1564, 12) & to_signed(-121922, 20)),
		std_logic_vector(to_signed(1566, 12) & to_signed(-120357, 20)),
		std_logic_vector(to_signed(1567, 12) & to_signed(-118791, 20)),
		std_logic_vector(to_signed(1568, 12) & to_signed(-117224, 20)),
		std_logic_vector(to_signed(1569, 12) & to_signed(-115656, 20)),
		std_logic_vector(to_signed(1570, 12) & to_signed(-114086, 20)),
		std_logic_vector(to_signed(1571, 12) & to_signed(-112516, 20)),
		std_logic_vector(to_signed(1572, 12) & to_signed(-110944, 20)),
		std_logic_vector(to_signed(1573, 12) & to_signed(-109372, 20)),
		std_logic_vector(to_signed(1574, 12) & to_signed(-107798, 20)),
		std_logic_vector(to_signed(1575, 12) & to_signed(-106224, 20)),
		std_logic_vector(to_signed(1576, 12) & to_signed(-104648, 20)),
		std_logic_vector(to_signed(1577, 12) & to_signed(-103071, 20)),
		std_logic_vector(to_signed(1578, 12) & to_signed(-101494, 20)),
		std_logic_vector(to_signed(1579, 12) & to_signed(-99915, 20)),
		std_logic_vector(to_signed(1580, 12) & to_signed(-98336, 20)),
		std_logic_vector(to_signed(1581, 12) & to_signed(-96755, 20)),
		std_logic_vector(to_signed(1582, 12) & to_signed(-95174, 20)),
		std_logic_vector(to_signed(1583, 12) & to_signed(-93592, 20)),
		std_logic_vector(to_signed(1584, 12) & to_signed(-92009, 20)),
		std_logic_vector(to_signed(1584, 12) & to_signed(-90425, 20)),
		std_logic_vector(to_signed(1585, 12) & to_signed(-88840, 20)),
		std_logic_vector(to_signed(1586, 12) & to_signed(-87254, 20)),
		std_logic_vector(to_signed(1587, 12) & to_signed(-85668, 20)),
		std_logic_vector(to_signed(1588, 12) & to_signed(-84081, 20)),
		std_logic_vector(to_signed(1588, 12) & to_signed(-82493, 20)),
		std_logic_vector(to_signed(1589, 12) & to_signed(-80904, 20)),
		std_logic_vector(to_signed(1590, 12) & to_signed(-79314, 20)),
		std_logic_vector(to_signed(1591, 12) & to_signed(-77724, 20)),
		std_logic_vector(to_signed(1591, 12) & to_signed(-76133, 20)),
		std_logic_vector(to_signed(1592, 12) & to_signed(-74541, 20)),
		std_logic_vector(to_signed(1593, 12) & to_signed(-72949, 20)),
		std_logic_vector(to_signed(1594, 12) & to_signed(-71355, 20)),
		std_logic_vector(to_signed(1594, 12) & to_signed(-69762, 20)),
		std_logic_vector(to_signed(1595, 12) & to_signed(-68167, 20)),
		std_logic_vector(to_signed(1595, 12) & to_signed(-66572, 20)),
		std_logic_vector(to_signed(1596, 12) & to_signed(-64976, 20)),
		std_logic_vector(to_signed(1597, 12) & to_signed(-63380, 20)),
		std_logic_vector(to_signed(1597, 12) & to_signed(-61783, 20)),
		std_logic_vector(to_signed(1598, 12) & to_signed(-60185, 20)),
		std_logic_vector(to_signed(1598, 12) & to_signed(-58587, 20)),
		std_logic_vector(to_signed(1599, 12) & to_signed(-56988, 20)),
		std_logic_vector(to_signed(1599, 12) & to_signed(-55389, 20)),
		std_logic_vector(to_signed(1600, 12) & to_signed(-53789, 20)),
		std_logic_vector(to_signed(1600, 12) & to_signed(-52189, 20)),
		std_logic_vector(to_signed(1601, 12) & to_signed(-50588, 20)),
		std_logic_vector(to_signed(1601, 12) & to_signed(-48987, 20)),
		std_logic_vector(to_signed(1602, 12) & to_signed(-47386, 20)),
		std_logic_vector(to_signed(1602, 12) & to_signed(-45783, 20)),
		std_logic_vector(to_signed(1603, 12) & to_signed(-44181, 20)),
		std_logic_vector(to_signed(1603, 12) & to_signed(-42578, 20)),
		std_logic_vector(to_signed(1604, 12) & to_signed(-40974, 20)),
		std_logic_vector(to_signed(1604, 12) & to_signed(-39371, 20)),
		std_logic_vector(to_signed(1604, 12) & to_signed(-37767, 20)),
		std_logic_vector(to_signed(1605, 12) & to_signed(-36162, 20)),
		std_logic_vector(to_signed(1605, 12) & to_signed(-34557, 20)),
		std_logic_vector(to_signed(1605, 12) & to_signed(-32952, 20)),
		std_logic_vector(to_signed(1606, 12) & to_signed(-31347, 20)),
		std_logic_vector(to_signed(1606, 12) & to_signed(-29741, 20)),
		std_logic_vector(to_signed(1606, 12) & to_signed(-28135, 20)),
		std_logic_vector(to_signed(1606, 12) & to_signed(-26529, 20)),
		std_logic_vector(to_signed(1607, 12) & to_signed(-24922, 20)),
		std_logic_vector(to_signed(1607, 12) & to_signed(-23315, 20)),
		std_logic_vector(to_signed(1607, 12) & to_signed(-21708, 20)),
		std_logic_vector(to_signed(1607, 12) & to_signed(-20101, 20)),
		std_logic_vector(to_signed(1607, 12) & to_signed(-18494, 20)),
		std_logic_vector(to_signed(1608, 12) & to_signed(-16886, 20)),
		std_logic_vector(to_signed(1608, 12) & to_signed(-15278, 20)),
		std_logic_vector(to_signed(1608, 12) & to_signed(-13671, 20)),
		std_logic_vector(to_signed(1608, 12) & to_signed(-12063, 20)),
		std_logic_vector(to_signed(1608, 12) & to_signed(-10454, 20)),
		std_logic_vector(to_signed(1608, 12) & to_signed(-8846, 20)),
		std_logic_vector(to_signed(1608, 12) & to_signed(-7238, 20)),
		std_logic_vector(to_signed(1608, 12) & to_signed(-5630, 20)),
		std_logic_vector(to_signed(1608, 12) & to_signed(-4021, 20)),
		std_logic_vector(to_signed(1608, 12) & to_signed(-2413, 20)),
		std_logic_vector(to_signed(1608, 12) & to_signed(-804, 20))
	);
	
	-- Signals
	signal TableAddrA	: std_logic_vector(log2ceil(TableSize_c)-1 downto 0);
	signal TableDataA	: std_logic_vector(TableWidth_c-1 downto 0);
	signal TableAddrB	: std_logic_vector(log2ceil(TableSize_c)-1 downto 0);
	signal TableDataB	: std_logic_vector(TableWidth_c-1 downto 0);
	
	
begin

	-- *** Calculation Unit ***
	i_calc_a : entity work.psi_fix_lin_approx_calc
		generic map (
			InFmt_g			=> InFmt_c,
			OutFmt_g		=> OutFmt_c,
			OffsFmt_g		=> OffsFmt_c,
			GradFmt_g		=> GradFmt_c,
			TableSize_g		=> TableSize_c
		)
		port map (
			-- Control Signals
			Clk			=> Clk,
			Rst			=> Rst,
			-- Input
			InVld		=> InVldA,
			InData		=> InDataA,
			-- Output
			OutVld		=> OutVldA,
			OutData		=> OutDataA,
			-- Table Interface
			TblAddr		=> TableAddrA,
			TblData		=> TableDataA
		);
	i_calc_b : entity work.psi_fix_lin_approx_calc
		generic map (
			InFmt_g			=> InFmt_c,
			OutFmt_g		=> OutFmt_c,
			OffsFmt_g		=> OffsFmt_c,
			GradFmt_g		=> GradFmt_c,
			TableSize_g		=> TableSize_c
		)
		port map (
			-- Control Signals
			Clk			=> Clk,
			Rst			=> Rst,
			-- Input
			InVld		=> InVldB,
			InData		=> InDataB,
			-- Output
			OutVld		=> OutVldB,
			OutData		=> OutDataB,
			-- Table Interface
			TblAddr		=> TableAddrB,
			TblData		=> TableDataB
		);		
	-- *** Table ***
	p_table : process(Clk)
	begin
		if rising_edge(Clk) then
			TableDataA <= Table_c(to_integer(unsigned(TableAddrA)));
			TableDataB <= Table_c(to_integer(unsigned(TableAddrB)));
		end if;
	end process;
	

end rtl;