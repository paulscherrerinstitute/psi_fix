------------------------------------------------------------------------------
--  Copyright (c) 2018 by Paul Scherrer Institute, Switzerland
--  All rights reserved.
------------------------------------------------------------------------------

------------------------------------------------------------------------------
-- Libraries
------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library work;
use work.psi_fix_pkg.all;
use work.psi_common_math_pkg.all;

------------------------------------------------------------------------------
-- Entity Declaration
------------------------------------------------------------------------------
entity psi_fix_lin_approx_gaussify20b is
  port(
    -- Control Signals
    Clk     : in  std_logic;
    Rst     : in  std_logic;
    -- Input
    InVld   : in  std_logic;
    InData  : in  std_logic_vector(20 - 1 downto 0); -- Format (1, 0, 19)
    -- Output
    OutVld  : out std_logic;
    OutData : out std_logic_vector(20 - 1 downto 0) -- Format (1, 0, 19)
  );
end entity;

------------------------------------------------------------------------------
-- Architecture Declaration
------------------------------------------------------------------------------
architecture rtl of psi_fix_lin_approx_gaussify20b is

  -- Constants
  constant InFmt_c      : PsiFixFmt_t := (1, 0, 19);
  constant OutFmt_c     : PsiFixFmt_t := (1, 0, 19);
  constant OffsFmt_c    : PsiFixFmt_t := (1, 0, 21);
  constant GradFmt_c    : PsiFixFmt_t := (0, 5, 9);
  constant TableSize_c  : integer     := 1024;
  constant TableWidth_c : integer     := 36;

  -- Table

  type Table_t is array (0 to TableSize_c - 1) of std_logic_vector(TableWidth_c - 1 downto 0);
  constant Table_c : Table_t := (
    std_logic_vector(to_signed(213, 14) & to_signed(854, 22)),
    std_logic_vector(to_signed(213, 14) & to_signed(2562, 22)),
    std_logic_vector(to_signed(213, 14) & to_signed(4269, 22)),
    std_logic_vector(to_signed(213, 14) & to_signed(5977, 22)),
    std_logic_vector(to_signed(213, 14) & to_signed(7685, 22)),
    std_logic_vector(to_signed(213, 14) & to_signed(9393, 22)),
    std_logic_vector(to_signed(213, 14) & to_signed(11101, 22)),
    std_logic_vector(to_signed(214, 14) & to_signed(12809, 22)),
    std_logic_vector(to_signed(214, 14) & to_signed(14517, 22)),
    std_logic_vector(to_signed(214, 14) & to_signed(16225, 22)),
    std_logic_vector(to_signed(214, 14) & to_signed(17934, 22)),
    std_logic_vector(to_signed(214, 14) & to_signed(19642, 22)),
    std_logic_vector(to_signed(214, 14) & to_signed(21350, 22)),
    std_logic_vector(to_signed(214, 14) & to_signed(23059, 22)),
    std_logic_vector(to_signed(214, 14) & to_signed(24768, 22)),
    std_logic_vector(to_signed(214, 14) & to_signed(26477, 22)),
    std_logic_vector(to_signed(214, 14) & to_signed(28186, 22)),
    std_logic_vector(to_signed(214, 14) & to_signed(29895, 22)),
    std_logic_vector(to_signed(214, 14) & to_signed(31605, 22)),
    std_logic_vector(to_signed(214, 14) & to_signed(33314, 22)),
    std_logic_vector(to_signed(214, 14) & to_signed(35024, 22)),
    std_logic_vector(to_signed(214, 14) & to_signed(36734, 22)),
    std_logic_vector(to_signed(214, 14) & to_signed(38444, 22)),
    std_logic_vector(to_signed(214, 14) & to_signed(40155, 22)),
    std_logic_vector(to_signed(214, 14) & to_signed(41865, 22)),
    std_logic_vector(to_signed(214, 14) & to_signed(43576, 22)),
    std_logic_vector(to_signed(214, 14) & to_signed(45288, 22)),
    std_logic_vector(to_signed(214, 14) & to_signed(46999, 22)),
    std_logic_vector(to_signed(214, 14) & to_signed(48711, 22)),
    std_logic_vector(to_signed(214, 14) & to_signed(50423, 22)),
    std_logic_vector(to_signed(214, 14) & to_signed(52135, 22)),
    std_logic_vector(to_signed(214, 14) & to_signed(53848, 22)),
    std_logic_vector(to_signed(214, 14) & to_signed(55561, 22)),
    std_logic_vector(to_signed(214, 14) & to_signed(57274, 22)),
    std_logic_vector(to_signed(214, 14) & to_signed(58988, 22)),
    std_logic_vector(to_signed(214, 14) & to_signed(60702, 22)),
    std_logic_vector(to_signed(214, 14) & to_signed(62416, 22)),
    std_logic_vector(to_signed(214, 14) & to_signed(64131, 22)),
    std_logic_vector(to_signed(214, 14) & to_signed(65846, 22)),
    std_logic_vector(to_signed(214, 14) & to_signed(67562, 22)),
    std_logic_vector(to_signed(215, 14) & to_signed(69278, 22)),
    std_logic_vector(to_signed(215, 14) & to_signed(70994, 22)),
    std_logic_vector(to_signed(215, 14) & to_signed(72711, 22)),
    std_logic_vector(to_signed(215, 14) & to_signed(74428, 22)),
    std_logic_vector(to_signed(215, 14) & to_signed(76146, 22)),
    std_logic_vector(to_signed(215, 14) & to_signed(77864, 22)),
    std_logic_vector(to_signed(215, 14) & to_signed(79583, 22)),
    std_logic_vector(to_signed(215, 14) & to_signed(81302, 22)),
    std_logic_vector(to_signed(215, 14) & to_signed(83022, 22)),
    std_logic_vector(to_signed(215, 14) & to_signed(84742, 22)),
    std_logic_vector(to_signed(215, 14) & to_signed(86462, 22)),
    std_logic_vector(to_signed(215, 14) & to_signed(88184, 22)),
    std_logic_vector(to_signed(215, 14) & to_signed(89905, 22)),
    std_logic_vector(to_signed(215, 14) & to_signed(91627, 22)),
    std_logic_vector(to_signed(215, 14) & to_signed(93350, 22)),
    std_logic_vector(to_signed(215, 14) & to_signed(95074, 22)),
    std_logic_vector(to_signed(216, 14) & to_signed(96797, 22)),
    std_logic_vector(to_signed(216, 14) & to_signed(98522, 22)),
    std_logic_vector(to_signed(216, 14) & to_signed(100247, 22)),
    std_logic_vector(to_signed(216, 14) & to_signed(101973, 22)),
    std_logic_vector(to_signed(216, 14) & to_signed(103699, 22)),
    std_logic_vector(to_signed(216, 14) & to_signed(105426, 22)),
    std_logic_vector(to_signed(216, 14) & to_signed(107154, 22)),
    std_logic_vector(to_signed(216, 14) & to_signed(108882, 22)),
    std_logic_vector(to_signed(216, 14) & to_signed(110611, 22)),
    std_logic_vector(to_signed(216, 14) & to_signed(112341, 22)),
    std_logic_vector(to_signed(216, 14) & to_signed(114071, 22)),
    std_logic_vector(to_signed(216, 14) & to_signed(115802, 22)),
    std_logic_vector(to_signed(217, 14) & to_signed(117534, 22)),
    std_logic_vector(to_signed(217, 14) & to_signed(119266, 22)),
    std_logic_vector(to_signed(217, 14) & to_signed(120999, 22)),
    std_logic_vector(to_signed(217, 14) & to_signed(122733, 22)),
    std_logic_vector(to_signed(217, 14) & to_signed(124468, 22)),
    std_logic_vector(to_signed(217, 14) & to_signed(126203, 22)),
    std_logic_vector(to_signed(217, 14) & to_signed(127940, 22)),
    std_logic_vector(to_signed(217, 14) & to_signed(129677, 22)),
    std_logic_vector(to_signed(217, 14) & to_signed(131414, 22)),
    std_logic_vector(to_signed(217, 14) & to_signed(133153, 22)),
    std_logic_vector(to_signed(217, 14) & to_signed(134892, 22)),
    std_logic_vector(to_signed(218, 14) & to_signed(136633, 22)),
    std_logic_vector(to_signed(218, 14) & to_signed(138374, 22)),
    std_logic_vector(to_signed(218, 14) & to_signed(140116, 22)),
    std_logic_vector(to_signed(218, 14) & to_signed(141859, 22)),
    std_logic_vector(to_signed(218, 14) & to_signed(143602, 22)),
    std_logic_vector(to_signed(218, 14) & to_signed(145347, 22)),
    std_logic_vector(to_signed(218, 14) & to_signed(147093, 22)),
    std_logic_vector(to_signed(218, 14) & to_signed(148839, 22)),
    std_logic_vector(to_signed(218, 14) & to_signed(150586, 22)),
    std_logic_vector(to_signed(219, 14) & to_signed(152335, 22)),
    std_logic_vector(to_signed(219, 14) & to_signed(154084, 22)),
    std_logic_vector(to_signed(219, 14) & to_signed(155834, 22)),
    std_logic_vector(to_signed(219, 14) & to_signed(157586, 22)),
    std_logic_vector(to_signed(219, 14) & to_signed(159338, 22)),
    std_logic_vector(to_signed(219, 14) & to_signed(161091, 22)),
    std_logic_vector(to_signed(219, 14) & to_signed(162845, 22)),
    std_logic_vector(to_signed(219, 14) & to_signed(164601, 22)),
    std_logic_vector(to_signed(220, 14) & to_signed(166357, 22)),
    std_logic_vector(to_signed(220, 14) & to_signed(168114, 22)),
    std_logic_vector(to_signed(220, 14) & to_signed(169873, 22)),
    std_logic_vector(to_signed(220, 14) & to_signed(171632, 22)),
    std_logic_vector(to_signed(220, 14) & to_signed(173393, 22)),
    std_logic_vector(to_signed(220, 14) & to_signed(175154, 22)),
    std_logic_vector(to_signed(220, 14) & to_signed(176917, 22)),
    std_logic_vector(to_signed(221, 14) & to_signed(178681, 22)),
    std_logic_vector(to_signed(221, 14) & to_signed(180446, 22)),
    std_logic_vector(to_signed(221, 14) & to_signed(182212, 22)),
    std_logic_vector(to_signed(221, 14) & to_signed(183980, 22)),
    std_logic_vector(to_signed(221, 14) & to_signed(185748, 22)),
    std_logic_vector(to_signed(221, 14) & to_signed(187518, 22)),
    std_logic_vector(to_signed(221, 14) & to_signed(189289, 22)),
    std_logic_vector(to_signed(222, 14) & to_signed(191061, 22)),
    std_logic_vector(to_signed(222, 14) & to_signed(192834, 22)),
    std_logic_vector(to_signed(222, 14) & to_signed(194609, 22)),
    std_logic_vector(to_signed(222, 14) & to_signed(196385, 22)),
    std_logic_vector(to_signed(222, 14) & to_signed(198162, 22)),
    std_logic_vector(to_signed(222, 14) & to_signed(199940, 22)),
    std_logic_vector(to_signed(223, 14) & to_signed(201720, 22)),
    std_logic_vector(to_signed(223, 14) & to_signed(203501, 22)),
    std_logic_vector(to_signed(223, 14) & to_signed(205284, 22)),
    std_logic_vector(to_signed(223, 14) & to_signed(207067, 22)),
    std_logic_vector(to_signed(223, 14) & to_signed(208852, 22)),
    std_logic_vector(to_signed(223, 14) & to_signed(210639, 22)),
    std_logic_vector(to_signed(224, 14) & to_signed(212426, 22)),
    std_logic_vector(to_signed(224, 14) & to_signed(214216, 22)),
    std_logic_vector(to_signed(224, 14) & to_signed(216006, 22)),
    std_logic_vector(to_signed(224, 14) & to_signed(217798, 22)),
    std_logic_vector(to_signed(224, 14) & to_signed(219592, 22)),
    std_logic_vector(to_signed(224, 14) & to_signed(221386, 22)),
    std_logic_vector(to_signed(225, 14) & to_signed(223183, 22)),
    std_logic_vector(to_signed(225, 14) & to_signed(224981, 22)),
    std_logic_vector(to_signed(225, 14) & to_signed(226780, 22)),
    std_logic_vector(to_signed(225, 14) & to_signed(228581, 22)),
    std_logic_vector(to_signed(225, 14) & to_signed(230383, 22)),
    std_logic_vector(to_signed(226, 14) & to_signed(232187, 22)),
    std_logic_vector(to_signed(226, 14) & to_signed(233992, 22)),
    std_logic_vector(to_signed(226, 14) & to_signed(235799, 22)),
    std_logic_vector(to_signed(226, 14) & to_signed(237608, 22)),
    std_logic_vector(to_signed(226, 14) & to_signed(239418, 22)),
    std_logic_vector(to_signed(227, 14) & to_signed(241230, 22)),
    std_logic_vector(to_signed(227, 14) & to_signed(243043, 22)),
    std_logic_vector(to_signed(227, 14) & to_signed(244858, 22)),
    std_logic_vector(to_signed(227, 14) & to_signed(246675, 22)),
    std_logic_vector(to_signed(227, 14) & to_signed(248493, 22)),
    std_logic_vector(to_signed(228, 14) & to_signed(250313, 22)),
    std_logic_vector(to_signed(228, 14) & to_signed(252135, 22)),
    std_logic_vector(to_signed(228, 14) & to_signed(253958, 22)),
    std_logic_vector(to_signed(228, 14) & to_signed(255783, 22)),
    std_logic_vector(to_signed(228, 14) & to_signed(257610, 22)),
    std_logic_vector(to_signed(229, 14) & to_signed(259439, 22)),
    std_logic_vector(to_signed(229, 14) & to_signed(261269, 22)),
    std_logic_vector(to_signed(229, 14) & to_signed(263101, 22)),
    std_logic_vector(to_signed(229, 14) & to_signed(264935, 22)),
    std_logic_vector(to_signed(230, 14) & to_signed(266771, 22)),
    std_logic_vector(to_signed(230, 14) & to_signed(268609, 22)),
    std_logic_vector(to_signed(230, 14) & to_signed(270448, 22)),
    std_logic_vector(to_signed(230, 14) & to_signed(272290, 22)),
    std_logic_vector(to_signed(231, 14) & to_signed(274133, 22)),
    std_logic_vector(to_signed(231, 14) & to_signed(275978, 22)),
    std_logic_vector(to_signed(231, 14) & to_signed(277825, 22)),
    std_logic_vector(to_signed(231, 14) & to_signed(279675, 22)),
    std_logic_vector(to_signed(232, 14) & to_signed(281526, 22)),
    std_logic_vector(to_signed(232, 14) & to_signed(283379, 22)),
    std_logic_vector(to_signed(232, 14) & to_signed(285234, 22)),
    std_logic_vector(to_signed(232, 14) & to_signed(287091, 22)),
    std_logic_vector(to_signed(233, 14) & to_signed(288950, 22)),
    std_logic_vector(to_signed(233, 14) & to_signed(290811, 22)),
    std_logic_vector(to_signed(233, 14) & to_signed(292674, 22)),
    std_logic_vector(to_signed(233, 14) & to_signed(294539, 22)),
    std_logic_vector(to_signed(234, 14) & to_signed(296407, 22)),
    std_logic_vector(to_signed(234, 14) & to_signed(298276, 22)),
    std_logic_vector(to_signed(234, 14) & to_signed(300148, 22)),
    std_logic_vector(to_signed(234, 14) & to_signed(302021, 22)),
    std_logic_vector(to_signed(235, 14) & to_signed(303897, 22)),
    std_logic_vector(to_signed(235, 14) & to_signed(305775, 22)),
    std_logic_vector(to_signed(235, 14) & to_signed(307656, 22)),
    std_logic_vector(to_signed(235, 14) & to_signed(309538, 22)),
    std_logic_vector(to_signed(236, 14) & to_signed(311423, 22)),
    std_logic_vector(to_signed(236, 14) & to_signed(313310, 22)),
    std_logic_vector(to_signed(236, 14) & to_signed(315199, 22)),
    std_logic_vector(to_signed(237, 14) & to_signed(317091, 22)),
    std_logic_vector(to_signed(237, 14) & to_signed(318985, 22)),
    std_logic_vector(to_signed(237, 14) & to_signed(320881, 22)),
    std_logic_vector(to_signed(237, 14) & to_signed(322780, 22)),
    std_logic_vector(to_signed(238, 14) & to_signed(324681, 22)),
    std_logic_vector(to_signed(238, 14) & to_signed(326585, 22)),
    std_logic_vector(to_signed(238, 14) & to_signed(328491, 22)),
    std_logic_vector(to_signed(239, 14) & to_signed(330399, 22)),
    std_logic_vector(to_signed(239, 14) & to_signed(332310, 22)),
    std_logic_vector(to_signed(239, 14) & to_signed(334223, 22)),
    std_logic_vector(to_signed(240, 14) & to_signed(336139, 22)),
    std_logic_vector(to_signed(240, 14) & to_signed(338057, 22)),
    std_logic_vector(to_signed(240, 14) & to_signed(339978, 22)),
    std_logic_vector(to_signed(241, 14) & to_signed(341902, 22)),
    std_logic_vector(to_signed(241, 14) & to_signed(343828, 22)),
    std_logic_vector(to_signed(241, 14) & to_signed(345756, 22)),
    std_logic_vector(to_signed(242, 14) & to_signed(347688, 22)),
    std_logic_vector(to_signed(242, 14) & to_signed(349622, 22)),
    std_logic_vector(to_signed(242, 14) & to_signed(351558, 22)),
    std_logic_vector(to_signed(243, 14) & to_signed(353498, 22)),
    std_logic_vector(to_signed(243, 14) & to_signed(355440, 22)),
    std_logic_vector(to_signed(243, 14) & to_signed(357384, 22)),
    std_logic_vector(to_signed(244, 14) & to_signed(359332, 22)),
    std_logic_vector(to_signed(244, 14) & to_signed(361282, 22)),
    std_logic_vector(to_signed(244, 14) & to_signed(363236, 22)),
    std_logic_vector(to_signed(245, 14) & to_signed(365192, 22)),
    std_logic_vector(to_signed(245, 14) & to_signed(367150, 22)),
    std_logic_vector(to_signed(245, 14) & to_signed(369112, 22)),
    std_logic_vector(to_signed(246, 14) & to_signed(371077, 22)),
    std_logic_vector(to_signed(246, 14) & to_signed(373045, 22)),
    std_logic_vector(to_signed(247, 14) & to_signed(375015, 22)),
    std_logic_vector(to_signed(247, 14) & to_signed(376989, 22)),
    std_logic_vector(to_signed(247, 14) & to_signed(378965, 22)),
    std_logic_vector(to_signed(248, 14) & to_signed(380945, 22)),
    std_logic_vector(to_signed(248, 14) & to_signed(382928, 22)),
    std_logic_vector(to_signed(248, 14) & to_signed(384913, 22)),
    std_logic_vector(to_signed(249, 14) & to_signed(386902, 22)),
    std_logic_vector(to_signed(249, 14) & to_signed(388894, 22)),
    std_logic_vector(to_signed(250, 14) & to_signed(390889, 22)),
    std_logic_vector(to_signed(250, 14) & to_signed(392888, 22)),
    std_logic_vector(to_signed(250, 14) & to_signed(394889, 22)),
    std_logic_vector(to_signed(251, 14) & to_signed(396894, 22)),
    std_logic_vector(to_signed(251, 14) & to_signed(398902, 22)),
    std_logic_vector(to_signed(252, 14) & to_signed(400914, 22)),
    std_logic_vector(to_signed(252, 14) & to_signed(402928, 22)),
    std_logic_vector(to_signed(252, 14) & to_signed(404946, 22)),
    std_logic_vector(to_signed(253, 14) & to_signed(406968, 22)),
    std_logic_vector(to_signed(253, 14) & to_signed(408993, 22)),
    std_logic_vector(to_signed(254, 14) & to_signed(411021, 22)),
    std_logic_vector(to_signed(254, 14) & to_signed(413053, 22)),
    std_logic_vector(to_signed(255, 14) & to_signed(415088, 22)),
    std_logic_vector(to_signed(255, 14) & to_signed(417127, 22)),
    std_logic_vector(to_signed(256, 14) & to_signed(419169, 22)),
    std_logic_vector(to_signed(256, 14) & to_signed(421215, 22)),
    std_logic_vector(to_signed(256, 14) & to_signed(423264, 22)),
    std_logic_vector(to_signed(257, 14) & to_signed(425318, 22)),
    std_logic_vector(to_signed(257, 14) & to_signed(427375, 22)),
    std_logic_vector(to_signed(258, 14) & to_signed(429435, 22)),
    std_logic_vector(to_signed(258, 14) & to_signed(431499, 22)),
    std_logic_vector(to_signed(259, 14) & to_signed(433567, 22)),
    std_logic_vector(to_signed(259, 14) & to_signed(435639, 22)),
    std_logic_vector(to_signed(260, 14) & to_signed(437715, 22)),
    std_logic_vector(to_signed(260, 14) & to_signed(439795, 22)),
    std_logic_vector(to_signed(261, 14) & to_signed(441878, 22)),
    std_logic_vector(to_signed(261, 14) & to_signed(443965, 22)),
    std_logic_vector(to_signed(262, 14) & to_signed(446057, 22)),
    std_logic_vector(to_signed(262, 14) & to_signed(448152, 22)),
    std_logic_vector(to_signed(263, 14) & to_signed(450252, 22)),
    std_logic_vector(to_signed(263, 14) & to_signed(452355, 22)),
    std_logic_vector(to_signed(264, 14) & to_signed(454463, 22)),
    std_logic_vector(to_signed(264, 14) & to_signed(456574, 22)),
    std_logic_vector(to_signed(265, 14) & to_signed(458690, 22)),
    std_logic_vector(to_signed(265, 14) & to_signed(460810, 22)),
    std_logic_vector(to_signed(266, 14) & to_signed(462935, 22)),
    std_logic_vector(to_signed(266, 14) & to_signed(465063, 22)),
    std_logic_vector(to_signed(267, 14) & to_signed(467196, 22)),
    std_logic_vector(to_signed(267, 14) & to_signed(469333, 22)),
    std_logic_vector(to_signed(268, 14) & to_signed(471475, 22)),
    std_logic_vector(to_signed(269, 14) & to_signed(473621, 22)),
    std_logic_vector(to_signed(269, 14) & to_signed(475772, 22)),
    std_logic_vector(to_signed(270, 14) & to_signed(477927, 22)),
    std_logic_vector(to_signed(270, 14) & to_signed(480087, 22)),
    std_logic_vector(to_signed(271, 14) & to_signed(482251, 22)),
    std_logic_vector(to_signed(271, 14) & to_signed(484420, 22)),
    std_logic_vector(to_signed(272, 14) & to_signed(486593, 22)),
    std_logic_vector(to_signed(273, 14) & to_signed(488772, 22)),
    std_logic_vector(to_signed(273, 14) & to_signed(490955, 22)),
    std_logic_vector(to_signed(274, 14) & to_signed(493143, 22)),
    std_logic_vector(to_signed(274, 14) & to_signed(495335, 22)),
    std_logic_vector(to_signed(275, 14) & to_signed(497533, 22)),
    std_logic_vector(to_signed(276, 14) & to_signed(499735, 22)),
    std_logic_vector(to_signed(276, 14) & to_signed(501943, 22)),
    std_logic_vector(to_signed(277, 14) & to_signed(504155, 22)),
    std_logic_vector(to_signed(278, 14) & to_signed(506373, 22)),
    std_logic_vector(to_signed(278, 14) & to_signed(508595, 22)),
    std_logic_vector(to_signed(279, 14) & to_signed(510823, 22)),
    std_logic_vector(to_signed(279, 14) & to_signed(513056, 22)),
    std_logic_vector(to_signed(280, 14) & to_signed(515295, 22)),
    std_logic_vector(to_signed(281, 14) & to_signed(517538, 22)),
    std_logic_vector(to_signed(281, 14) & to_signed(519787, 22)),
    std_logic_vector(to_signed(282, 14) & to_signed(522041, 22)),
    std_logic_vector(to_signed(283, 14) & to_signed(524301, 22)),
    std_logic_vector(to_signed(283, 14) & to_signed(526566, 22)),
    std_logic_vector(to_signed(284, 14) & to_signed(528837, 22)),
    std_logic_vector(to_signed(285, 14) & to_signed(531113, 22)),
    std_logic_vector(to_signed(286, 14) & to_signed(533395, 22)),
    std_logic_vector(to_signed(286, 14) & to_signed(535683, 22)),
    std_logic_vector(to_signed(287, 14) & to_signed(537976, 22)),
    std_logic_vector(to_signed(288, 14) & to_signed(540276, 22)),
    std_logic_vector(to_signed(289, 14) & to_signed(542581, 22)),
    std_logic_vector(to_signed(289, 14) & to_signed(544892, 22)),
    std_logic_vector(to_signed(290, 14) & to_signed(547209, 22)),
    std_logic_vector(to_signed(291, 14) & to_signed(549532, 22)),
    std_logic_vector(to_signed(292, 14) & to_signed(551861, 22)),
    std_logic_vector(to_signed(292, 14) & to_signed(554196, 22)),
    std_logic_vector(to_signed(293, 14) & to_signed(556538, 22)),
    std_logic_vector(to_signed(294, 14) & to_signed(558885, 22)),
    std_logic_vector(to_signed(295, 14) & to_signed(561239, 22)),
    std_logic_vector(to_signed(295, 14) & to_signed(563600, 22)),
    std_logic_vector(to_signed(296, 14) & to_signed(565967, 22)),
    std_logic_vector(to_signed(297, 14) & to_signed(568340, 22)),
    std_logic_vector(to_signed(298, 14) & to_signed(570720, 22)),
    std_logic_vector(to_signed(299, 14) & to_signed(573107, 22)),
    std_logic_vector(to_signed(300, 14) & to_signed(575500, 22)),
    std_logic_vector(to_signed(300, 14) & to_signed(577900, 22)),
    std_logic_vector(to_signed(301, 14) & to_signed(580307, 22)),
    std_logic_vector(to_signed(302, 14) & to_signed(582721, 22)),
    std_logic_vector(to_signed(303, 14) & to_signed(585141, 22)),
    std_logic_vector(to_signed(304, 14) & to_signed(587569, 22)),
    std_logic_vector(to_signed(305, 14) & to_signed(590004, 22)),
    std_logic_vector(to_signed(306, 14) & to_signed(592446, 22)),
    std_logic_vector(to_signed(307, 14) & to_signed(594895, 22)),
    std_logic_vector(to_signed(308, 14) & to_signed(597352, 22)),
    std_logic_vector(to_signed(308, 14) & to_signed(599816, 22)),
    std_logic_vector(to_signed(309, 14) & to_signed(602287, 22)),
    std_logic_vector(to_signed(310, 14) & to_signed(604767, 22)),
    std_logic_vector(to_signed(311, 14) & to_signed(607253, 22)),
    std_logic_vector(to_signed(312, 14) & to_signed(609748, 22)),
    std_logic_vector(to_signed(313, 14) & to_signed(612250, 22)),
    std_logic_vector(to_signed(314, 14) & to_signed(614760, 22)),
    std_logic_vector(to_signed(315, 14) & to_signed(617278, 22)),
    std_logic_vector(to_signed(316, 14) & to_signed(619804, 22)),
    std_logic_vector(to_signed(317, 14) & to_signed(622338, 22)),
    std_logic_vector(to_signed(318, 14) & to_signed(624880, 22)),
    std_logic_vector(to_signed(319, 14) & to_signed(627431, 22)),
    std_logic_vector(to_signed(320, 14) & to_signed(629990, 22)),
    std_logic_vector(to_signed(321, 14) & to_signed(632558, 22)),
    std_logic_vector(to_signed(323, 14) & to_signed(635134, 22)),
    std_logic_vector(to_signed(324, 14) & to_signed(637718, 22)),
    std_logic_vector(to_signed(325, 14) & to_signed(640312, 22)),
    std_logic_vector(to_signed(326, 14) & to_signed(642914, 22)),
    std_logic_vector(to_signed(327, 14) & to_signed(645525, 22)),
    std_logic_vector(to_signed(328, 14) & to_signed(648146, 22)),
    std_logic_vector(to_signed(329, 14) & to_signed(650775, 22)),
    std_logic_vector(to_signed(330, 14) & to_signed(653414, 22)),
    std_logic_vector(to_signed(332, 14) & to_signed(656062, 22)),
    std_logic_vector(to_signed(333, 14) & to_signed(658719, 22)),
    std_logic_vector(to_signed(334, 14) & to_signed(661386, 22)),
    std_logic_vector(to_signed(335, 14) & to_signed(664063, 22)),
    std_logic_vector(to_signed(336, 14) & to_signed(666749, 22)),
    std_logic_vector(to_signed(338, 14) & to_signed(669446, 22)),
    std_logic_vector(to_signed(339, 14) & to_signed(672152, 22)),
    std_logic_vector(to_signed(340, 14) & to_signed(674869, 22)),
    std_logic_vector(to_signed(341, 14) & to_signed(677595, 22)),
    std_logic_vector(to_signed(343, 14) & to_signed(680332, 22)),
    std_logic_vector(to_signed(344, 14) & to_signed(683080, 22)),
    std_logic_vector(to_signed(345, 14) & to_signed(685838, 22)),
    std_logic_vector(to_signed(347, 14) & to_signed(688607, 22)),
    std_logic_vector(to_signed(348, 14) & to_signed(691386, 22)),
    std_logic_vector(to_signed(350, 14) & to_signed(694177, 22)),
    std_logic_vector(to_signed(351, 14) & to_signed(696979, 22)),
    std_logic_vector(to_signed(352, 14) & to_signed(699792, 22)),
    std_logic_vector(to_signed(354, 14) & to_signed(702616, 22)),
    std_logic_vector(to_signed(355, 14) & to_signed(705452, 22)),
    std_logic_vector(to_signed(357, 14) & to_signed(708299, 22)),
    std_logic_vector(to_signed(358, 14) & to_signed(711159, 22)),
    std_logic_vector(to_signed(360, 14) & to_signed(714030, 22)),
    std_logic_vector(to_signed(361, 14) & to_signed(716913, 22)),
    std_logic_vector(to_signed(363, 14) & to_signed(719809, 22)),
    std_logic_vector(to_signed(364, 14) & to_signed(722717, 22)),
    std_logic_vector(to_signed(366, 14) & to_signed(725637, 22)),
    std_logic_vector(to_signed(367, 14) & to_signed(728571, 22)),
    std_logic_vector(to_signed(369, 14) & to_signed(731517, 22)),
    std_logic_vector(to_signed(371, 14) & to_signed(734476, 22)),
    std_logic_vector(to_signed(372, 14) & to_signed(737449, 22)),
    std_logic_vector(to_signed(374, 14) & to_signed(740435, 22)),
    std_logic_vector(to_signed(376, 14) & to_signed(743434, 22)),
    std_logic_vector(to_signed(378, 14) & to_signed(746447, 22)),
    std_logic_vector(to_signed(379, 14) & to_signed(749474, 22)),
    std_logic_vector(to_signed(381, 14) & to_signed(752515, 22)),
    std_logic_vector(to_signed(383, 14) & to_signed(755571, 22)),
    std_logic_vector(to_signed(385, 14) & to_signed(758641, 22)),
    std_logic_vector(to_signed(387, 14) & to_signed(761726, 22)),
    std_logic_vector(to_signed(388, 14) & to_signed(764825, 22)),
    std_logic_vector(to_signed(390, 14) & to_signed(767940, 22)),
    std_logic_vector(to_signed(392, 14) & to_signed(771070, 22)),
    std_logic_vector(to_signed(394, 14) & to_signed(774216, 22)),
    std_logic_vector(to_signed(396, 14) & to_signed(777377, 22)),
    std_logic_vector(to_signed(398, 14) & to_signed(780555, 22)),
    std_logic_vector(to_signed(400, 14) & to_signed(783748, 22)),
    std_logic_vector(to_signed(402, 14) & to_signed(786958, 22)),
    std_logic_vector(to_signed(404, 14) & to_signed(790185, 22)),
    std_logic_vector(to_signed(407, 14) & to_signed(793428, 22)),
    std_logic_vector(to_signed(409, 14) & to_signed(796689, 22)),
    std_logic_vector(to_signed(411, 14) & to_signed(799967, 22)),
    std_logic_vector(to_signed(413, 14) & to_signed(803263, 22)),
    std_logic_vector(to_signed(415, 14) & to_signed(806577, 22)),
    std_logic_vector(to_signed(418, 14) & to_signed(809909, 22)),
    std_logic_vector(to_signed(420, 14) & to_signed(813260, 22)),
    std_logic_vector(to_signed(422, 14) & to_signed(816629, 22)),
    std_logic_vector(to_signed(425, 14) & to_signed(820018, 22)),
    std_logic_vector(to_signed(427, 14) & to_signed(823425, 22)),
    std_logic_vector(to_signed(430, 14) & to_signed(826853, 22)),
    std_logic_vector(to_signed(432, 14) & to_signed(830300, 22)),
    std_logic_vector(to_signed(435, 14) & to_signed(833768, 22)),
    std_logic_vector(to_signed(437, 14) & to_signed(837257, 22)),
    std_logic_vector(to_signed(440, 14) & to_signed(840766, 22)),
    std_logic_vector(to_signed(443, 14) & to_signed(844297, 22)),
    std_logic_vector(to_signed(445, 14) & to_signed(847849, 22)),
    std_logic_vector(to_signed(448, 14) & to_signed(851424, 22)),
    std_logic_vector(to_signed(451, 14) & to_signed(855021, 22)),
    std_logic_vector(to_signed(454, 14) & to_signed(858640, 22)),
    std_logic_vector(to_signed(457, 14) & to_signed(862283, 22)),
    std_logic_vector(to_signed(460, 14) & to_signed(865949, 22)),
    std_logic_vector(to_signed(463, 14) & to_signed(869640, 22)),
    std_logic_vector(to_signed(466, 14) & to_signed(873355, 22)),
    std_logic_vector(to_signed(469, 14) & to_signed(877094, 22)),
    std_logic_vector(to_signed(472, 14) & to_signed(880859, 22)),
    std_logic_vector(to_signed(475, 14) & to_signed(884650, 22)),
    std_logic_vector(to_signed(479, 14) & to_signed(888466, 22)),
    std_logic_vector(to_signed(482, 14) & to_signed(892310, 22)),
    std_logic_vector(to_signed(486, 14) & to_signed(896180, 22)),
    std_logic_vector(to_signed(489, 14) & to_signed(900079, 22)),
    std_logic_vector(to_signed(493, 14) & to_signed(904005, 22)),
    std_logic_vector(to_signed(496, 14) & to_signed(907960, 22)),
    std_logic_vector(to_signed(500, 14) & to_signed(911945, 22)),
    std_logic_vector(to_signed(504, 14) & to_signed(915959, 22)),
    std_logic_vector(to_signed(508, 14) & to_signed(920004, 22)),
    std_logic_vector(to_signed(511, 14) & to_signed(924080, 22)),
    std_logic_vector(to_signed(515, 14) & to_signed(928187, 22)),
    std_logic_vector(to_signed(520, 14) & to_signed(932327, 22)),
    std_logic_vector(to_signed(524, 14) & to_signed(936500, 22)),
    std_logic_vector(to_signed(528, 14) & to_signed(940706, 22)),
    std_logic_vector(to_signed(532, 14) & to_signed(944947, 22)),
    std_logic_vector(to_signed(537, 14) & to_signed(949222, 22)),
    std_logic_vector(to_signed(541, 14) & to_signed(953534, 22)),
    std_logic_vector(to_signed(546, 14) & to_signed(957882, 22)),
    std_logic_vector(to_signed(551, 14) & to_signed(962268, 22)),
    std_logic_vector(to_signed(555, 14) & to_signed(966691, 22)),
    std_logic_vector(to_signed(560, 14) & to_signed(971154, 22)),
    std_logic_vector(to_signed(565, 14) & to_signed(975657, 22)),
    std_logic_vector(to_signed(571, 14) & to_signed(980200, 22)),
    std_logic_vector(to_signed(576, 14) & to_signed(984786, 22)),
    std_logic_vector(to_signed(581, 14) & to_signed(989414, 22)),
    std_logic_vector(to_signed(587, 14) & to_signed(994086, 22)),
    std_logic_vector(to_signed(592, 14) & to_signed(998803, 22)),
    std_logic_vector(to_signed(598, 14) & to_signed(1003565, 22)),
    std_logic_vector(to_signed(604, 14) & to_signed(1008375, 22)),
    std_logic_vector(to_signed(610, 14) & to_signed(1013233, 22)),
    std_logic_vector(to_signed(617, 14) & to_signed(1018140, 22)),
    std_logic_vector(to_signed(623, 14) & to_signed(1023098, 22)),
    std_logic_vector(to_signed(630, 14) & to_signed(1028109, 22)),
    std_logic_vector(to_signed(636, 14) & to_signed(1033172, 22)),
    std_logic_vector(to_signed(643, 14) & to_signed(1038290, 22)),
    std_logic_vector(to_signed(650, 14) & to_signed(1043465, 22)),
    std_logic_vector(to_signed(658, 14) & to_signed(1048697, 22)),
    std_logic_vector(to_signed(665, 14) & to_signed(1053989, 22)),
    std_logic_vector(to_signed(673, 14) & to_signed(1059342, 22)),
    std_logic_vector(to_signed(681, 14) & to_signed(1064758, 22)),
    std_logic_vector(to_signed(689, 14) & to_signed(1070238, 22)),
    std_logic_vector(to_signed(698, 14) & to_signed(1075785, 22)),
    std_logic_vector(to_signed(706, 14) & to_signed(1081400, 22)),
    std_logic_vector(to_signed(715, 14) & to_signed(1087087, 22)),
    std_logic_vector(to_signed(725, 14) & to_signed(1092846, 22)),
    std_logic_vector(to_signed(734, 14) & to_signed(1098680, 22)),
    std_logic_vector(to_signed(744, 14) & to_signed(1104592, 22)),
    std_logic_vector(to_signed(754, 14) & to_signed(1110584, 22)),
    std_logic_vector(to_signed(765, 14) & to_signed(1116658, 22)),
    std_logic_vector(to_signed(775, 14) & to_signed(1122818, 22)),
    std_logic_vector(to_signed(787, 14) & to_signed(1129067, 22)),
    std_logic_vector(to_signed(798, 14) & to_signed(1135407, 22)),
    std_logic_vector(to_signed(810, 14) & to_signed(1141842, 22)),
    std_logic_vector(to_signed(823, 14) & to_signed(1148375, 22)),
    std_logic_vector(to_signed(836, 14) & to_signed(1155010, 22)),
    std_logic_vector(to_signed(849, 14) & to_signed(1161751, 22)),
    std_logic_vector(to_signed(863, 14) & to_signed(1168602, 22)),
    std_logic_vector(to_signed(878, 14) & to_signed(1175566, 22)),
    std_logic_vector(to_signed(893, 14) & to_signed(1182650, 22)),
    std_logic_vector(to_signed(909, 14) & to_signed(1189857, 22)),
    std_logic_vector(to_signed(925, 14) & to_signed(1197192, 22)),
    std_logic_vector(to_signed(942, 14) & to_signed(1204662, 22)),
    std_logic_vector(to_signed(960, 14) & to_signed(1212273, 22)),
    std_logic_vector(to_signed(979, 14) & to_signed(1220029, 22)),
    std_logic_vector(to_signed(999, 14) & to_signed(1227939, 22)),
    std_logic_vector(to_signed(1019, 14) & to_signed(1236009, 22)),
    std_logic_vector(to_signed(1041, 14) & to_signed(1244248, 22)),
    std_logic_vector(to_signed(1063, 14) & to_signed(1252663, 22)),
    std_logic_vector(to_signed(1087, 14) & to_signed(1261264, 22)),
    std_logic_vector(to_signed(1112, 14) & to_signed(1270060, 22)),
    std_logic_vector(to_signed(1138, 14) & to_signed(1279061, 22)),
    std_logic_vector(to_signed(1166, 14) & to_signed(1288280, 22)),
    std_logic_vector(to_signed(1196, 14) & to_signed(1297729, 22)),
    std_logic_vector(to_signed(1227, 14) & to_signed(1307421, 22)),
    std_logic_vector(to_signed(1260, 14) & to_signed(1317372, 22)),
    std_logic_vector(to_signed(1296, 14) & to_signed(1327596, 22)),
    std_logic_vector(to_signed(1333, 14) & to_signed(1338113, 22)),
    std_logic_vector(to_signed(1374, 14) & to_signed(1348942, 22)),
    std_logic_vector(to_signed(1417, 14) & to_signed(1360104, 22)),
    std_logic_vector(to_signed(1463, 14) & to_signed(1371625, 22)),
    std_logic_vector(to_signed(1513, 14) & to_signed(1383531, 22)),
    std_logic_vector(to_signed(1567, 14) & to_signed(1395853, 22)),
    std_logic_vector(to_signed(1626, 14) & to_signed(1408624, 22)),
    std_logic_vector(to_signed(1689, 14) & to_signed(1421884, 22)),
    std_logic_vector(to_signed(1759, 14) & to_signed(1435677, 22)),
    std_logic_vector(to_signed(1835, 14) & to_signed(1450052, 22)),
    std_logic_vector(to_signed(1919, 14) & to_signed(1465069, 22)),
    std_logic_vector(to_signed(2012, 14) & to_signed(1480794, 22)),
    std_logic_vector(to_signed(2116, 14) & to_signed(1497308, 22)),
    std_logic_vector(to_signed(2233, 14) & to_signed(1514702, 22)),
    std_logic_vector(to_signed(2364, 14) & to_signed(1533090, 22)),
    std_logic_vector(to_signed(2514, 14) & to_signed(1552605, 22)),
    std_logic_vector(to_signed(2687, 14) & to_signed(1573413, 22)),
    std_logic_vector(to_signed(2889, 14) & to_signed(1595719, 22)),
    std_logic_vector(to_signed(3127, 14) & to_signed(1619782, 22)),
    std_logic_vector(to_signed(3412, 14) & to_signed(1645938, 22)),
    std_logic_vector(to_signed(3761, 14) & to_signed(1674633, 22)),
    std_logic_vector(to_signed(4199, 14) & to_signed(1706474, 22)),
    std_logic_vector(to_signed(4764, 14) & to_signed(1742328, 22)),
    std_logic_vector(to_signed(5526, 14) & to_signed(1783488, 22)),
    std_logic_vector(to_signed(6609, 14) & to_signed(1832027, 22)),
    std_logic_vector(to_signed(8285, 14) & to_signed(1891606, 22)),
    std_logic_vector(to_signed(11256, 14) & to_signed(1969772, 22)),
    std_logic_vector(to_signed(10294, 14) & to_signed(2055974, 22)),
    std_logic_vector(to_signed(10294, 14) & to_signed(-2055974, 22)),
    std_logic_vector(to_signed(11256, 14) & to_signed(-1969772, 22)),
    std_logic_vector(to_signed(8285, 14) & to_signed(-1891606, 22)),
    std_logic_vector(to_signed(6609, 14) & to_signed(-1832027, 22)),
    std_logic_vector(to_signed(5526, 14) & to_signed(-1783488, 22)),
    std_logic_vector(to_signed(4764, 14) & to_signed(-1742328, 22)),
    std_logic_vector(to_signed(4199, 14) & to_signed(-1706474, 22)),
    std_logic_vector(to_signed(3761, 14) & to_signed(-1674633, 22)),
    std_logic_vector(to_signed(3412, 14) & to_signed(-1645938, 22)),
    std_logic_vector(to_signed(3127, 14) & to_signed(-1619782, 22)),
    std_logic_vector(to_signed(2889, 14) & to_signed(-1595719, 22)),
    std_logic_vector(to_signed(2687, 14) & to_signed(-1573413, 22)),
    std_logic_vector(to_signed(2514, 14) & to_signed(-1552605, 22)),
    std_logic_vector(to_signed(2364, 14) & to_signed(-1533090, 22)),
    std_logic_vector(to_signed(2233, 14) & to_signed(-1514702, 22)),
    std_logic_vector(to_signed(2116, 14) & to_signed(-1497308, 22)),
    std_logic_vector(to_signed(2012, 14) & to_signed(-1480794, 22)),
    std_logic_vector(to_signed(1919, 14) & to_signed(-1465069, 22)),
    std_logic_vector(to_signed(1835, 14) & to_signed(-1450052, 22)),
    std_logic_vector(to_signed(1759, 14) & to_signed(-1435677, 22)),
    std_logic_vector(to_signed(1689, 14) & to_signed(-1421884, 22)),
    std_logic_vector(to_signed(1626, 14) & to_signed(-1408624, 22)),
    std_logic_vector(to_signed(1567, 14) & to_signed(-1395853, 22)),
    std_logic_vector(to_signed(1513, 14) & to_signed(-1383531, 22)),
    std_logic_vector(to_signed(1463, 14) & to_signed(-1371625, 22)),
    std_logic_vector(to_signed(1417, 14) & to_signed(-1360104, 22)),
    std_logic_vector(to_signed(1374, 14) & to_signed(-1348942, 22)),
    std_logic_vector(to_signed(1333, 14) & to_signed(-1338113, 22)),
    std_logic_vector(to_signed(1296, 14) & to_signed(-1327596, 22)),
    std_logic_vector(to_signed(1260, 14) & to_signed(-1317372, 22)),
    std_logic_vector(to_signed(1227, 14) & to_signed(-1307421, 22)),
    std_logic_vector(to_signed(1196, 14) & to_signed(-1297729, 22)),
    std_logic_vector(to_signed(1166, 14) & to_signed(-1288280, 22)),
    std_logic_vector(to_signed(1138, 14) & to_signed(-1279061, 22)),
    std_logic_vector(to_signed(1112, 14) & to_signed(-1270060, 22)),
    std_logic_vector(to_signed(1087, 14) & to_signed(-1261264, 22)),
    std_logic_vector(to_signed(1063, 14) & to_signed(-1252663, 22)),
    std_logic_vector(to_signed(1041, 14) & to_signed(-1244248, 22)),
    std_logic_vector(to_signed(1019, 14) & to_signed(-1236009, 22)),
    std_logic_vector(to_signed(999, 14) & to_signed(-1227939, 22)),
    std_logic_vector(to_signed(979, 14) & to_signed(-1220029, 22)),
    std_logic_vector(to_signed(960, 14) & to_signed(-1212273, 22)),
    std_logic_vector(to_signed(942, 14) & to_signed(-1204662, 22)),
    std_logic_vector(to_signed(925, 14) & to_signed(-1197192, 22)),
    std_logic_vector(to_signed(909, 14) & to_signed(-1189857, 22)),
    std_logic_vector(to_signed(893, 14) & to_signed(-1182650, 22)),
    std_logic_vector(to_signed(878, 14) & to_signed(-1175566, 22)),
    std_logic_vector(to_signed(863, 14) & to_signed(-1168602, 22)),
    std_logic_vector(to_signed(849, 14) & to_signed(-1161751, 22)),
    std_logic_vector(to_signed(836, 14) & to_signed(-1155010, 22)),
    std_logic_vector(to_signed(823, 14) & to_signed(-1148375, 22)),
    std_logic_vector(to_signed(810, 14) & to_signed(-1141842, 22)),
    std_logic_vector(to_signed(798, 14) & to_signed(-1135407, 22)),
    std_logic_vector(to_signed(787, 14) & to_signed(-1129067, 22)),
    std_logic_vector(to_signed(775, 14) & to_signed(-1122818, 22)),
    std_logic_vector(to_signed(765, 14) & to_signed(-1116658, 22)),
    std_logic_vector(to_signed(754, 14) & to_signed(-1110584, 22)),
    std_logic_vector(to_signed(744, 14) & to_signed(-1104592, 22)),
    std_logic_vector(to_signed(734, 14) & to_signed(-1098680, 22)),
    std_logic_vector(to_signed(725, 14) & to_signed(-1092846, 22)),
    std_logic_vector(to_signed(715, 14) & to_signed(-1087087, 22)),
    std_logic_vector(to_signed(706, 14) & to_signed(-1081400, 22)),
    std_logic_vector(to_signed(698, 14) & to_signed(-1075785, 22)),
    std_logic_vector(to_signed(689, 14) & to_signed(-1070238, 22)),
    std_logic_vector(to_signed(681, 14) & to_signed(-1064758, 22)),
    std_logic_vector(to_signed(673, 14) & to_signed(-1059342, 22)),
    std_logic_vector(to_signed(665, 14) & to_signed(-1053989, 22)),
    std_logic_vector(to_signed(658, 14) & to_signed(-1048697, 22)),
    std_logic_vector(to_signed(650, 14) & to_signed(-1043465, 22)),
    std_logic_vector(to_signed(643, 14) & to_signed(-1038290, 22)),
    std_logic_vector(to_signed(636, 14) & to_signed(-1033172, 22)),
    std_logic_vector(to_signed(630, 14) & to_signed(-1028109, 22)),
    std_logic_vector(to_signed(623, 14) & to_signed(-1023098, 22)),
    std_logic_vector(to_signed(617, 14) & to_signed(-1018140, 22)),
    std_logic_vector(to_signed(610, 14) & to_signed(-1013233, 22)),
    std_logic_vector(to_signed(604, 14) & to_signed(-1008375, 22)),
    std_logic_vector(to_signed(598, 14) & to_signed(-1003565, 22)),
    std_logic_vector(to_signed(592, 14) & to_signed(-998803, 22)),
    std_logic_vector(to_signed(587, 14) & to_signed(-994086, 22)),
    std_logic_vector(to_signed(581, 14) & to_signed(-989414, 22)),
    std_logic_vector(to_signed(576, 14) & to_signed(-984786, 22)),
    std_logic_vector(to_signed(571, 14) & to_signed(-980200, 22)),
    std_logic_vector(to_signed(565, 14) & to_signed(-975657, 22)),
    std_logic_vector(to_signed(560, 14) & to_signed(-971154, 22)),
    std_logic_vector(to_signed(555, 14) & to_signed(-966691, 22)),
    std_logic_vector(to_signed(551, 14) & to_signed(-962268, 22)),
    std_logic_vector(to_signed(546, 14) & to_signed(-957882, 22)),
    std_logic_vector(to_signed(541, 14) & to_signed(-953534, 22)),
    std_logic_vector(to_signed(537, 14) & to_signed(-949222, 22)),
    std_logic_vector(to_signed(532, 14) & to_signed(-944947, 22)),
    std_logic_vector(to_signed(528, 14) & to_signed(-940706, 22)),
    std_logic_vector(to_signed(524, 14) & to_signed(-936500, 22)),
    std_logic_vector(to_signed(520, 14) & to_signed(-932327, 22)),
    std_logic_vector(to_signed(515, 14) & to_signed(-928187, 22)),
    std_logic_vector(to_signed(511, 14) & to_signed(-924080, 22)),
    std_logic_vector(to_signed(508, 14) & to_signed(-920004, 22)),
    std_logic_vector(to_signed(504, 14) & to_signed(-915959, 22)),
    std_logic_vector(to_signed(500, 14) & to_signed(-911945, 22)),
    std_logic_vector(to_signed(496, 14) & to_signed(-907960, 22)),
    std_logic_vector(to_signed(493, 14) & to_signed(-904005, 22)),
    std_logic_vector(to_signed(489, 14) & to_signed(-900079, 22)),
    std_logic_vector(to_signed(486, 14) & to_signed(-896180, 22)),
    std_logic_vector(to_signed(482, 14) & to_signed(-892310, 22)),
    std_logic_vector(to_signed(479, 14) & to_signed(-888466, 22)),
    std_logic_vector(to_signed(475, 14) & to_signed(-884650, 22)),
    std_logic_vector(to_signed(472, 14) & to_signed(-880859, 22)),
    std_logic_vector(to_signed(469, 14) & to_signed(-877094, 22)),
    std_logic_vector(to_signed(466, 14) & to_signed(-873355, 22)),
    std_logic_vector(to_signed(463, 14) & to_signed(-869640, 22)),
    std_logic_vector(to_signed(460, 14) & to_signed(-865949, 22)),
    std_logic_vector(to_signed(457, 14) & to_signed(-862283, 22)),
    std_logic_vector(to_signed(454, 14) & to_signed(-858640, 22)),
    std_logic_vector(to_signed(451, 14) & to_signed(-855021, 22)),
    std_logic_vector(to_signed(448, 14) & to_signed(-851424, 22)),
    std_logic_vector(to_signed(445, 14) & to_signed(-847849, 22)),
    std_logic_vector(to_signed(443, 14) & to_signed(-844297, 22)),
    std_logic_vector(to_signed(440, 14) & to_signed(-840766, 22)),
    std_logic_vector(to_signed(437, 14) & to_signed(-837257, 22)),
    std_logic_vector(to_signed(435, 14) & to_signed(-833768, 22)),
    std_logic_vector(to_signed(432, 14) & to_signed(-830300, 22)),
    std_logic_vector(to_signed(430, 14) & to_signed(-826853, 22)),
    std_logic_vector(to_signed(427, 14) & to_signed(-823425, 22)),
    std_logic_vector(to_signed(425, 14) & to_signed(-820018, 22)),
    std_logic_vector(to_signed(422, 14) & to_signed(-816629, 22)),
    std_logic_vector(to_signed(420, 14) & to_signed(-813260, 22)),
    std_logic_vector(to_signed(418, 14) & to_signed(-809909, 22)),
    std_logic_vector(to_signed(415, 14) & to_signed(-806577, 22)),
    std_logic_vector(to_signed(413, 14) & to_signed(-803263, 22)),
    std_logic_vector(to_signed(411, 14) & to_signed(-799967, 22)),
    std_logic_vector(to_signed(409, 14) & to_signed(-796689, 22)),
    std_logic_vector(to_signed(407, 14) & to_signed(-793428, 22)),
    std_logic_vector(to_signed(404, 14) & to_signed(-790185, 22)),
    std_logic_vector(to_signed(402, 14) & to_signed(-786958, 22)),
    std_logic_vector(to_signed(400, 14) & to_signed(-783748, 22)),
    std_logic_vector(to_signed(398, 14) & to_signed(-780555, 22)),
    std_logic_vector(to_signed(396, 14) & to_signed(-777377, 22)),
    std_logic_vector(to_signed(394, 14) & to_signed(-774216, 22)),
    std_logic_vector(to_signed(392, 14) & to_signed(-771070, 22)),
    std_logic_vector(to_signed(390, 14) & to_signed(-767940, 22)),
    std_logic_vector(to_signed(388, 14) & to_signed(-764825, 22)),
    std_logic_vector(to_signed(387, 14) & to_signed(-761726, 22)),
    std_logic_vector(to_signed(385, 14) & to_signed(-758641, 22)),
    std_logic_vector(to_signed(383, 14) & to_signed(-755571, 22)),
    std_logic_vector(to_signed(381, 14) & to_signed(-752515, 22)),
    std_logic_vector(to_signed(379, 14) & to_signed(-749474, 22)),
    std_logic_vector(to_signed(378, 14) & to_signed(-746447, 22)),
    std_logic_vector(to_signed(376, 14) & to_signed(-743434, 22)),
    std_logic_vector(to_signed(374, 14) & to_signed(-740435, 22)),
    std_logic_vector(to_signed(372, 14) & to_signed(-737449, 22)),
    std_logic_vector(to_signed(371, 14) & to_signed(-734476, 22)),
    std_logic_vector(to_signed(369, 14) & to_signed(-731517, 22)),
    std_logic_vector(to_signed(367, 14) & to_signed(-728571, 22)),
    std_logic_vector(to_signed(366, 14) & to_signed(-725637, 22)),
    std_logic_vector(to_signed(364, 14) & to_signed(-722717, 22)),
    std_logic_vector(to_signed(363, 14) & to_signed(-719809, 22)),
    std_logic_vector(to_signed(361, 14) & to_signed(-716913, 22)),
    std_logic_vector(to_signed(360, 14) & to_signed(-714030, 22)),
    std_logic_vector(to_signed(358, 14) & to_signed(-711159, 22)),
    std_logic_vector(to_signed(357, 14) & to_signed(-708299, 22)),
    std_logic_vector(to_signed(355, 14) & to_signed(-705452, 22)),
    std_logic_vector(to_signed(354, 14) & to_signed(-702616, 22)),
    std_logic_vector(to_signed(352, 14) & to_signed(-699792, 22)),
    std_logic_vector(to_signed(351, 14) & to_signed(-696979, 22)),
    std_logic_vector(to_signed(350, 14) & to_signed(-694177, 22)),
    std_logic_vector(to_signed(348, 14) & to_signed(-691386, 22)),
    std_logic_vector(to_signed(347, 14) & to_signed(-688607, 22)),
    std_logic_vector(to_signed(345, 14) & to_signed(-685838, 22)),
    std_logic_vector(to_signed(344, 14) & to_signed(-683080, 22)),
    std_logic_vector(to_signed(343, 14) & to_signed(-680332, 22)),
    std_logic_vector(to_signed(341, 14) & to_signed(-677595, 22)),
    std_logic_vector(to_signed(340, 14) & to_signed(-674869, 22)),
    std_logic_vector(to_signed(339, 14) & to_signed(-672152, 22)),
    std_logic_vector(to_signed(338, 14) & to_signed(-669446, 22)),
    std_logic_vector(to_signed(336, 14) & to_signed(-666749, 22)),
    std_logic_vector(to_signed(335, 14) & to_signed(-664063, 22)),
    std_logic_vector(to_signed(334, 14) & to_signed(-661386, 22)),
    std_logic_vector(to_signed(333, 14) & to_signed(-658719, 22)),
    std_logic_vector(to_signed(332, 14) & to_signed(-656062, 22)),
    std_logic_vector(to_signed(330, 14) & to_signed(-653414, 22)),
    std_logic_vector(to_signed(329, 14) & to_signed(-650775, 22)),
    std_logic_vector(to_signed(328, 14) & to_signed(-648146, 22)),
    std_logic_vector(to_signed(327, 14) & to_signed(-645525, 22)),
    std_logic_vector(to_signed(326, 14) & to_signed(-642914, 22)),
    std_logic_vector(to_signed(325, 14) & to_signed(-640312, 22)),
    std_logic_vector(to_signed(324, 14) & to_signed(-637718, 22)),
    std_logic_vector(to_signed(323, 14) & to_signed(-635134, 22)),
    std_logic_vector(to_signed(321, 14) & to_signed(-632558, 22)),
    std_logic_vector(to_signed(320, 14) & to_signed(-629990, 22)),
    std_logic_vector(to_signed(319, 14) & to_signed(-627431, 22)),
    std_logic_vector(to_signed(318, 14) & to_signed(-624880, 22)),
    std_logic_vector(to_signed(317, 14) & to_signed(-622338, 22)),
    std_logic_vector(to_signed(316, 14) & to_signed(-619804, 22)),
    std_logic_vector(to_signed(315, 14) & to_signed(-617278, 22)),
    std_logic_vector(to_signed(314, 14) & to_signed(-614760, 22)),
    std_logic_vector(to_signed(313, 14) & to_signed(-612250, 22)),
    std_logic_vector(to_signed(312, 14) & to_signed(-609748, 22)),
    std_logic_vector(to_signed(311, 14) & to_signed(-607253, 22)),
    std_logic_vector(to_signed(310, 14) & to_signed(-604767, 22)),
    std_logic_vector(to_signed(309, 14) & to_signed(-602287, 22)),
    std_logic_vector(to_signed(308, 14) & to_signed(-599816, 22)),
    std_logic_vector(to_signed(308, 14) & to_signed(-597352, 22)),
    std_logic_vector(to_signed(307, 14) & to_signed(-594895, 22)),
    std_logic_vector(to_signed(306, 14) & to_signed(-592446, 22)),
    std_logic_vector(to_signed(305, 14) & to_signed(-590004, 22)),
    std_logic_vector(to_signed(304, 14) & to_signed(-587569, 22)),
    std_logic_vector(to_signed(303, 14) & to_signed(-585141, 22)),
    std_logic_vector(to_signed(302, 14) & to_signed(-582721, 22)),
    std_logic_vector(to_signed(301, 14) & to_signed(-580307, 22)),
    std_logic_vector(to_signed(300, 14) & to_signed(-577900, 22)),
    std_logic_vector(to_signed(300, 14) & to_signed(-575500, 22)),
    std_logic_vector(to_signed(299, 14) & to_signed(-573107, 22)),
    std_logic_vector(to_signed(298, 14) & to_signed(-570720, 22)),
    std_logic_vector(to_signed(297, 14) & to_signed(-568340, 22)),
    std_logic_vector(to_signed(296, 14) & to_signed(-565967, 22)),
    std_logic_vector(to_signed(295, 14) & to_signed(-563600, 22)),
    std_logic_vector(to_signed(295, 14) & to_signed(-561239, 22)),
    std_logic_vector(to_signed(294, 14) & to_signed(-558885, 22)),
    std_logic_vector(to_signed(293, 14) & to_signed(-556538, 22)),
    std_logic_vector(to_signed(292, 14) & to_signed(-554196, 22)),
    std_logic_vector(to_signed(292, 14) & to_signed(-551861, 22)),
    std_logic_vector(to_signed(291, 14) & to_signed(-549532, 22)),
    std_logic_vector(to_signed(290, 14) & to_signed(-547209, 22)),
    std_logic_vector(to_signed(289, 14) & to_signed(-544892, 22)),
    std_logic_vector(to_signed(289, 14) & to_signed(-542581, 22)),
    std_logic_vector(to_signed(288, 14) & to_signed(-540276, 22)),
    std_logic_vector(to_signed(287, 14) & to_signed(-537976, 22)),
    std_logic_vector(to_signed(286, 14) & to_signed(-535683, 22)),
    std_logic_vector(to_signed(286, 14) & to_signed(-533395, 22)),
    std_logic_vector(to_signed(285, 14) & to_signed(-531113, 22)),
    std_logic_vector(to_signed(284, 14) & to_signed(-528837, 22)),
    std_logic_vector(to_signed(283, 14) & to_signed(-526566, 22)),
    std_logic_vector(to_signed(283, 14) & to_signed(-524301, 22)),
    std_logic_vector(to_signed(282, 14) & to_signed(-522041, 22)),
    std_logic_vector(to_signed(281, 14) & to_signed(-519787, 22)),
    std_logic_vector(to_signed(281, 14) & to_signed(-517538, 22)),
    std_logic_vector(to_signed(280, 14) & to_signed(-515295, 22)),
    std_logic_vector(to_signed(279, 14) & to_signed(-513056, 22)),
    std_logic_vector(to_signed(279, 14) & to_signed(-510823, 22)),
    std_logic_vector(to_signed(278, 14) & to_signed(-508595, 22)),
    std_logic_vector(to_signed(278, 14) & to_signed(-506373, 22)),
    std_logic_vector(to_signed(277, 14) & to_signed(-504155, 22)),
    std_logic_vector(to_signed(276, 14) & to_signed(-501943, 22)),
    std_logic_vector(to_signed(276, 14) & to_signed(-499735, 22)),
    std_logic_vector(to_signed(275, 14) & to_signed(-497533, 22)),
    std_logic_vector(to_signed(274, 14) & to_signed(-495335, 22)),
    std_logic_vector(to_signed(274, 14) & to_signed(-493143, 22)),
    std_logic_vector(to_signed(273, 14) & to_signed(-490955, 22)),
    std_logic_vector(to_signed(273, 14) & to_signed(-488772, 22)),
    std_logic_vector(to_signed(272, 14) & to_signed(-486593, 22)),
    std_logic_vector(to_signed(271, 14) & to_signed(-484420, 22)),
    std_logic_vector(to_signed(271, 14) & to_signed(-482251, 22)),
    std_logic_vector(to_signed(270, 14) & to_signed(-480087, 22)),
    std_logic_vector(to_signed(270, 14) & to_signed(-477927, 22)),
    std_logic_vector(to_signed(269, 14) & to_signed(-475772, 22)),
    std_logic_vector(to_signed(269, 14) & to_signed(-473621, 22)),
    std_logic_vector(to_signed(268, 14) & to_signed(-471475, 22)),
    std_logic_vector(to_signed(267, 14) & to_signed(-469333, 22)),
    std_logic_vector(to_signed(267, 14) & to_signed(-467196, 22)),
    std_logic_vector(to_signed(266, 14) & to_signed(-465063, 22)),
    std_logic_vector(to_signed(266, 14) & to_signed(-462935, 22)),
    std_logic_vector(to_signed(265, 14) & to_signed(-460810, 22)),
    std_logic_vector(to_signed(265, 14) & to_signed(-458690, 22)),
    std_logic_vector(to_signed(264, 14) & to_signed(-456574, 22)),
    std_logic_vector(to_signed(264, 14) & to_signed(-454463, 22)),
    std_logic_vector(to_signed(263, 14) & to_signed(-452355, 22)),
    std_logic_vector(to_signed(263, 14) & to_signed(-450252, 22)),
    std_logic_vector(to_signed(262, 14) & to_signed(-448152, 22)),
    std_logic_vector(to_signed(262, 14) & to_signed(-446057, 22)),
    std_logic_vector(to_signed(261, 14) & to_signed(-443965, 22)),
    std_logic_vector(to_signed(261, 14) & to_signed(-441878, 22)),
    std_logic_vector(to_signed(260, 14) & to_signed(-439795, 22)),
    std_logic_vector(to_signed(260, 14) & to_signed(-437715, 22)),
    std_logic_vector(to_signed(259, 14) & to_signed(-435639, 22)),
    std_logic_vector(to_signed(259, 14) & to_signed(-433567, 22)),
    std_logic_vector(to_signed(258, 14) & to_signed(-431499, 22)),
    std_logic_vector(to_signed(258, 14) & to_signed(-429435, 22)),
    std_logic_vector(to_signed(257, 14) & to_signed(-427375, 22)),
    std_logic_vector(to_signed(257, 14) & to_signed(-425318, 22)),
    std_logic_vector(to_signed(256, 14) & to_signed(-423264, 22)),
    std_logic_vector(to_signed(256, 14) & to_signed(-421215, 22)),
    std_logic_vector(to_signed(256, 14) & to_signed(-419169, 22)),
    std_logic_vector(to_signed(255, 14) & to_signed(-417127, 22)),
    std_logic_vector(to_signed(255, 14) & to_signed(-415088, 22)),
    std_logic_vector(to_signed(254, 14) & to_signed(-413053, 22)),
    std_logic_vector(to_signed(254, 14) & to_signed(-411021, 22)),
    std_logic_vector(to_signed(253, 14) & to_signed(-408993, 22)),
    std_logic_vector(to_signed(253, 14) & to_signed(-406968, 22)),
    std_logic_vector(to_signed(252, 14) & to_signed(-404946, 22)),
    std_logic_vector(to_signed(252, 14) & to_signed(-402928, 22)),
    std_logic_vector(to_signed(252, 14) & to_signed(-400914, 22)),
    std_logic_vector(to_signed(251, 14) & to_signed(-398902, 22)),
    std_logic_vector(to_signed(251, 14) & to_signed(-396894, 22)),
    std_logic_vector(to_signed(250, 14) & to_signed(-394889, 22)),
    std_logic_vector(to_signed(250, 14) & to_signed(-392888, 22)),
    std_logic_vector(to_signed(250, 14) & to_signed(-390889, 22)),
    std_logic_vector(to_signed(249, 14) & to_signed(-388894, 22)),
    std_logic_vector(to_signed(249, 14) & to_signed(-386902, 22)),
    std_logic_vector(to_signed(248, 14) & to_signed(-384913, 22)),
    std_logic_vector(to_signed(248, 14) & to_signed(-382928, 22)),
    std_logic_vector(to_signed(248, 14) & to_signed(-380945, 22)),
    std_logic_vector(to_signed(247, 14) & to_signed(-378965, 22)),
    std_logic_vector(to_signed(247, 14) & to_signed(-376989, 22)),
    std_logic_vector(to_signed(247, 14) & to_signed(-375015, 22)),
    std_logic_vector(to_signed(246, 14) & to_signed(-373045, 22)),
    std_logic_vector(to_signed(246, 14) & to_signed(-371077, 22)),
    std_logic_vector(to_signed(245, 14) & to_signed(-369112, 22)),
    std_logic_vector(to_signed(245, 14) & to_signed(-367150, 22)),
    std_logic_vector(to_signed(245, 14) & to_signed(-365192, 22)),
    std_logic_vector(to_signed(244, 14) & to_signed(-363236, 22)),
    std_logic_vector(to_signed(244, 14) & to_signed(-361282, 22)),
    std_logic_vector(to_signed(244, 14) & to_signed(-359332, 22)),
    std_logic_vector(to_signed(243, 14) & to_signed(-357384, 22)),
    std_logic_vector(to_signed(243, 14) & to_signed(-355440, 22)),
    std_logic_vector(to_signed(243, 14) & to_signed(-353498, 22)),
    std_logic_vector(to_signed(242, 14) & to_signed(-351558, 22)),
    std_logic_vector(to_signed(242, 14) & to_signed(-349622, 22)),
    std_logic_vector(to_signed(242, 14) & to_signed(-347688, 22)),
    std_logic_vector(to_signed(241, 14) & to_signed(-345756, 22)),
    std_logic_vector(to_signed(241, 14) & to_signed(-343828, 22)),
    std_logic_vector(to_signed(241, 14) & to_signed(-341902, 22)),
    std_logic_vector(to_signed(240, 14) & to_signed(-339978, 22)),
    std_logic_vector(to_signed(240, 14) & to_signed(-338057, 22)),
    std_logic_vector(to_signed(240, 14) & to_signed(-336139, 22)),
    std_logic_vector(to_signed(239, 14) & to_signed(-334223, 22)),
    std_logic_vector(to_signed(239, 14) & to_signed(-332310, 22)),
    std_logic_vector(to_signed(239, 14) & to_signed(-330399, 22)),
    std_logic_vector(to_signed(238, 14) & to_signed(-328491, 22)),
    std_logic_vector(to_signed(238, 14) & to_signed(-326585, 22)),
    std_logic_vector(to_signed(238, 14) & to_signed(-324681, 22)),
    std_logic_vector(to_signed(237, 14) & to_signed(-322780, 22)),
    std_logic_vector(to_signed(237, 14) & to_signed(-320881, 22)),
    std_logic_vector(to_signed(237, 14) & to_signed(-318985, 22)),
    std_logic_vector(to_signed(237, 14) & to_signed(-317091, 22)),
    std_logic_vector(to_signed(236, 14) & to_signed(-315199, 22)),
    std_logic_vector(to_signed(236, 14) & to_signed(-313310, 22)),
    std_logic_vector(to_signed(236, 14) & to_signed(-311423, 22)),
    std_logic_vector(to_signed(235, 14) & to_signed(-309538, 22)),
    std_logic_vector(to_signed(235, 14) & to_signed(-307656, 22)),
    std_logic_vector(to_signed(235, 14) & to_signed(-305775, 22)),
    std_logic_vector(to_signed(235, 14) & to_signed(-303897, 22)),
    std_logic_vector(to_signed(234, 14) & to_signed(-302021, 22)),
    std_logic_vector(to_signed(234, 14) & to_signed(-300148, 22)),
    std_logic_vector(to_signed(234, 14) & to_signed(-298276, 22)),
    std_logic_vector(to_signed(234, 14) & to_signed(-296407, 22)),
    std_logic_vector(to_signed(233, 14) & to_signed(-294539, 22)),
    std_logic_vector(to_signed(233, 14) & to_signed(-292674, 22)),
    std_logic_vector(to_signed(233, 14) & to_signed(-290811, 22)),
    std_logic_vector(to_signed(233, 14) & to_signed(-288950, 22)),
    std_logic_vector(to_signed(232, 14) & to_signed(-287091, 22)),
    std_logic_vector(to_signed(232, 14) & to_signed(-285234, 22)),
    std_logic_vector(to_signed(232, 14) & to_signed(-283379, 22)),
    std_logic_vector(to_signed(232, 14) & to_signed(-281526, 22)),
    std_logic_vector(to_signed(231, 14) & to_signed(-279675, 22)),
    std_logic_vector(to_signed(231, 14) & to_signed(-277825, 22)),
    std_logic_vector(to_signed(231, 14) & to_signed(-275978, 22)),
    std_logic_vector(to_signed(231, 14) & to_signed(-274133, 22)),
    std_logic_vector(to_signed(230, 14) & to_signed(-272290, 22)),
    std_logic_vector(to_signed(230, 14) & to_signed(-270448, 22)),
    std_logic_vector(to_signed(230, 14) & to_signed(-268609, 22)),
    std_logic_vector(to_signed(230, 14) & to_signed(-266771, 22)),
    std_logic_vector(to_signed(229, 14) & to_signed(-264935, 22)),
    std_logic_vector(to_signed(229, 14) & to_signed(-263101, 22)),
    std_logic_vector(to_signed(229, 14) & to_signed(-261269, 22)),
    std_logic_vector(to_signed(229, 14) & to_signed(-259439, 22)),
    std_logic_vector(to_signed(228, 14) & to_signed(-257610, 22)),
    std_logic_vector(to_signed(228, 14) & to_signed(-255783, 22)),
    std_logic_vector(to_signed(228, 14) & to_signed(-253958, 22)),
    std_logic_vector(to_signed(228, 14) & to_signed(-252135, 22)),
    std_logic_vector(to_signed(228, 14) & to_signed(-250313, 22)),
    std_logic_vector(to_signed(227, 14) & to_signed(-248493, 22)),
    std_logic_vector(to_signed(227, 14) & to_signed(-246675, 22)),
    std_logic_vector(to_signed(227, 14) & to_signed(-244858, 22)),
    std_logic_vector(to_signed(227, 14) & to_signed(-243043, 22)),
    std_logic_vector(to_signed(227, 14) & to_signed(-241230, 22)),
    std_logic_vector(to_signed(226, 14) & to_signed(-239418, 22)),
    std_logic_vector(to_signed(226, 14) & to_signed(-237608, 22)),
    std_logic_vector(to_signed(226, 14) & to_signed(-235799, 22)),
    std_logic_vector(to_signed(226, 14) & to_signed(-233992, 22)),
    std_logic_vector(to_signed(226, 14) & to_signed(-232187, 22)),
    std_logic_vector(to_signed(225, 14) & to_signed(-230383, 22)),
    std_logic_vector(to_signed(225, 14) & to_signed(-228581, 22)),
    std_logic_vector(to_signed(225, 14) & to_signed(-226780, 22)),
    std_logic_vector(to_signed(225, 14) & to_signed(-224981, 22)),
    std_logic_vector(to_signed(225, 14) & to_signed(-223183, 22)),
    std_logic_vector(to_signed(224, 14) & to_signed(-221386, 22)),
    std_logic_vector(to_signed(224, 14) & to_signed(-219592, 22)),
    std_logic_vector(to_signed(224, 14) & to_signed(-217798, 22)),
    std_logic_vector(to_signed(224, 14) & to_signed(-216006, 22)),
    std_logic_vector(to_signed(224, 14) & to_signed(-214216, 22)),
    std_logic_vector(to_signed(224, 14) & to_signed(-212426, 22)),
    std_logic_vector(to_signed(223, 14) & to_signed(-210639, 22)),
    std_logic_vector(to_signed(223, 14) & to_signed(-208852, 22)),
    std_logic_vector(to_signed(223, 14) & to_signed(-207067, 22)),
    std_logic_vector(to_signed(223, 14) & to_signed(-205284, 22)),
    std_logic_vector(to_signed(223, 14) & to_signed(-203501, 22)),
    std_logic_vector(to_signed(223, 14) & to_signed(-201720, 22)),
    std_logic_vector(to_signed(222, 14) & to_signed(-199940, 22)),
    std_logic_vector(to_signed(222, 14) & to_signed(-198162, 22)),
    std_logic_vector(to_signed(222, 14) & to_signed(-196385, 22)),
    std_logic_vector(to_signed(222, 14) & to_signed(-194609, 22)),
    std_logic_vector(to_signed(222, 14) & to_signed(-192834, 22)),
    std_logic_vector(to_signed(222, 14) & to_signed(-191061, 22)),
    std_logic_vector(to_signed(221, 14) & to_signed(-189289, 22)),
    std_logic_vector(to_signed(221, 14) & to_signed(-187518, 22)),
    std_logic_vector(to_signed(221, 14) & to_signed(-185748, 22)),
    std_logic_vector(to_signed(221, 14) & to_signed(-183980, 22)),
    std_logic_vector(to_signed(221, 14) & to_signed(-182212, 22)),
    std_logic_vector(to_signed(221, 14) & to_signed(-180446, 22)),
    std_logic_vector(to_signed(221, 14) & to_signed(-178681, 22)),
    std_logic_vector(to_signed(220, 14) & to_signed(-176917, 22)),
    std_logic_vector(to_signed(220, 14) & to_signed(-175154, 22)),
    std_logic_vector(to_signed(220, 14) & to_signed(-173393, 22)),
    std_logic_vector(to_signed(220, 14) & to_signed(-171632, 22)),
    std_logic_vector(to_signed(220, 14) & to_signed(-169873, 22)),
    std_logic_vector(to_signed(220, 14) & to_signed(-168114, 22)),
    std_logic_vector(to_signed(220, 14) & to_signed(-166357, 22)),
    std_logic_vector(to_signed(219, 14) & to_signed(-164601, 22)),
    std_logic_vector(to_signed(219, 14) & to_signed(-162845, 22)),
    std_logic_vector(to_signed(219, 14) & to_signed(-161091, 22)),
    std_logic_vector(to_signed(219, 14) & to_signed(-159338, 22)),
    std_logic_vector(to_signed(219, 14) & to_signed(-157586, 22)),
    std_logic_vector(to_signed(219, 14) & to_signed(-155834, 22)),
    std_logic_vector(to_signed(219, 14) & to_signed(-154084, 22)),
    std_logic_vector(to_signed(219, 14) & to_signed(-152335, 22)),
    std_logic_vector(to_signed(218, 14) & to_signed(-150586, 22)),
    std_logic_vector(to_signed(218, 14) & to_signed(-148839, 22)),
    std_logic_vector(to_signed(218, 14) & to_signed(-147093, 22)),
    std_logic_vector(to_signed(218, 14) & to_signed(-145347, 22)),
    std_logic_vector(to_signed(218, 14) & to_signed(-143602, 22)),
    std_logic_vector(to_signed(218, 14) & to_signed(-141859, 22)),
    std_logic_vector(to_signed(218, 14) & to_signed(-140116, 22)),
    std_logic_vector(to_signed(218, 14) & to_signed(-138374, 22)),
    std_logic_vector(to_signed(218, 14) & to_signed(-136633, 22)),
    std_logic_vector(to_signed(217, 14) & to_signed(-134892, 22)),
    std_logic_vector(to_signed(217, 14) & to_signed(-133153, 22)),
    std_logic_vector(to_signed(217, 14) & to_signed(-131414, 22)),
    std_logic_vector(to_signed(217, 14) & to_signed(-129677, 22)),
    std_logic_vector(to_signed(217, 14) & to_signed(-127940, 22)),
    std_logic_vector(to_signed(217, 14) & to_signed(-126203, 22)),
    std_logic_vector(to_signed(217, 14) & to_signed(-124468, 22)),
    std_logic_vector(to_signed(217, 14) & to_signed(-122733, 22)),
    std_logic_vector(to_signed(217, 14) & to_signed(-120999, 22)),
    std_logic_vector(to_signed(217, 14) & to_signed(-119266, 22)),
    std_logic_vector(to_signed(217, 14) & to_signed(-117534, 22)),
    std_logic_vector(to_signed(216, 14) & to_signed(-115802, 22)),
    std_logic_vector(to_signed(216, 14) & to_signed(-114071, 22)),
    std_logic_vector(to_signed(216, 14) & to_signed(-112341, 22)),
    std_logic_vector(to_signed(216, 14) & to_signed(-110611, 22)),
    std_logic_vector(to_signed(216, 14) & to_signed(-108882, 22)),
    std_logic_vector(to_signed(216, 14) & to_signed(-107154, 22)),
    std_logic_vector(to_signed(216, 14) & to_signed(-105426, 22)),
    std_logic_vector(to_signed(216, 14) & to_signed(-103699, 22)),
    std_logic_vector(to_signed(216, 14) & to_signed(-101973, 22)),
    std_logic_vector(to_signed(216, 14) & to_signed(-100247, 22)),
    std_logic_vector(to_signed(216, 14) & to_signed(-98522, 22)),
    std_logic_vector(to_signed(216, 14) & to_signed(-96797, 22)),
    std_logic_vector(to_signed(215, 14) & to_signed(-95074, 22)),
    std_logic_vector(to_signed(215, 14) & to_signed(-93350, 22)),
    std_logic_vector(to_signed(215, 14) & to_signed(-91627, 22)),
    std_logic_vector(to_signed(215, 14) & to_signed(-89905, 22)),
    std_logic_vector(to_signed(215, 14) & to_signed(-88184, 22)),
    std_logic_vector(to_signed(215, 14) & to_signed(-86462, 22)),
    std_logic_vector(to_signed(215, 14) & to_signed(-84742, 22)),
    std_logic_vector(to_signed(215, 14) & to_signed(-83022, 22)),
    std_logic_vector(to_signed(215, 14) & to_signed(-81302, 22)),
    std_logic_vector(to_signed(215, 14) & to_signed(-79583, 22)),
    std_logic_vector(to_signed(215, 14) & to_signed(-77864, 22)),
    std_logic_vector(to_signed(215, 14) & to_signed(-76146, 22)),
    std_logic_vector(to_signed(215, 14) & to_signed(-74428, 22)),
    std_logic_vector(to_signed(215, 14) & to_signed(-72711, 22)),
    std_logic_vector(to_signed(215, 14) & to_signed(-70994, 22)),
    std_logic_vector(to_signed(215, 14) & to_signed(-69278, 22)),
    std_logic_vector(to_signed(214, 14) & to_signed(-67562, 22)),
    std_logic_vector(to_signed(214, 14) & to_signed(-65846, 22)),
    std_logic_vector(to_signed(214, 14) & to_signed(-64131, 22)),
    std_logic_vector(to_signed(214, 14) & to_signed(-62416, 22)),
    std_logic_vector(to_signed(214, 14) & to_signed(-60702, 22)),
    std_logic_vector(to_signed(214, 14) & to_signed(-58988, 22)),
    std_logic_vector(to_signed(214, 14) & to_signed(-57274, 22)),
    std_logic_vector(to_signed(214, 14) & to_signed(-55561, 22)),
    std_logic_vector(to_signed(214, 14) & to_signed(-53848, 22)),
    std_logic_vector(to_signed(214, 14) & to_signed(-52135, 22)),
    std_logic_vector(to_signed(214, 14) & to_signed(-50423, 22)),
    std_logic_vector(to_signed(214, 14) & to_signed(-48711, 22)),
    std_logic_vector(to_signed(214, 14) & to_signed(-46999, 22)),
    std_logic_vector(to_signed(214, 14) & to_signed(-45288, 22)),
    std_logic_vector(to_signed(214, 14) & to_signed(-43576, 22)),
    std_logic_vector(to_signed(214, 14) & to_signed(-41865, 22)),
    std_logic_vector(to_signed(214, 14) & to_signed(-40155, 22)),
    std_logic_vector(to_signed(214, 14) & to_signed(-38444, 22)),
    std_logic_vector(to_signed(214, 14) & to_signed(-36734, 22)),
    std_logic_vector(to_signed(214, 14) & to_signed(-35024, 22)),
    std_logic_vector(to_signed(214, 14) & to_signed(-33314, 22)),
    std_logic_vector(to_signed(214, 14) & to_signed(-31605, 22)),
    std_logic_vector(to_signed(214, 14) & to_signed(-29895, 22)),
    std_logic_vector(to_signed(214, 14) & to_signed(-28186, 22)),
    std_logic_vector(to_signed(214, 14) & to_signed(-26477, 22)),
    std_logic_vector(to_signed(214, 14) & to_signed(-24768, 22)),
    std_logic_vector(to_signed(214, 14) & to_signed(-23059, 22)),
    std_logic_vector(to_signed(214, 14) & to_signed(-21350, 22)),
    std_logic_vector(to_signed(214, 14) & to_signed(-19642, 22)),
    std_logic_vector(to_signed(214, 14) & to_signed(-17934, 22)),
    std_logic_vector(to_signed(214, 14) & to_signed(-16225, 22)),
    std_logic_vector(to_signed(214, 14) & to_signed(-14517, 22)),
    std_logic_vector(to_signed(214, 14) & to_signed(-12809, 22)),
    std_logic_vector(to_signed(213, 14) & to_signed(-11101, 22)),
    std_logic_vector(to_signed(213, 14) & to_signed(-9393, 22)),
    std_logic_vector(to_signed(213, 14) & to_signed(-7685, 22)),
    std_logic_vector(to_signed(213, 14) & to_signed(-5977, 22)),
    std_logic_vector(to_signed(213, 14) & to_signed(-4269, 22)),
    std_logic_vector(to_signed(213, 14) & to_signed(-2562, 22)),
    std_logic_vector(to_signed(213, 14) & to_signed(-854, 22))
  );

  -- Signals
  signal TableAddr : std_logic_vector(log2ceil(TableSize_c) - 1 downto 0);
  signal TableData : std_logic_vector(TableWidth_c - 1 downto 0);

begin

  -- *** Calculation Unit ***
  i_calc : entity work.psi_fix_lin_approx_calc
    generic map(
      InFmt_g     => InFmt_c,
      OutFmt_g    => OutFmt_c,
      OffsFmt_g   => OffsFmt_c,
      GradFmt_g   => GradFmt_c,
      TableSize_g => TableSize_c
    )
    port map(
      -- Control Signals
      Clk     => Clk,
      Rst     => Rst,
      -- Input
      InVld   => InVld,
      InData  => InData,
      -- Output
      OutVld  => OutVld,
      OutData => OutData,
      -- Table Interface
      TblAddr => TableAddr,
      TblData => TableData
    );

  -- *** Table ***
  p_table : process(Clk)
  begin
    if rising_edge(Clk) then
      TableData <= Table_c(to_integer(unsigned(TableAddr)));
    end if;
  end process;

end architecture;
