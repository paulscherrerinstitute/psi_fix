------------------------------------------------------------------------------
--  Copyright (c) 2021 by Paul Scherrer Institute, Switzerland
--  All rights reserved.
--  Authors: Benoit Stef
------------------------------------------------------------------------------

------------------------------------------------------------------------------
-- Description
------------------------------------------------------------------------------
-- This block allows generating triggers out of several "analog" input signals
-- with fixed point format and several external triggers
-- The number of trigger generated is also extendable - quite specific though
-- intetntion to be used with multi stream DAQ
------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

use work.psi_common_math_pkg.all;
use work.psi_fix_pkg.all;
use work.psi_common_array_pkg.all;

--@formatter:off
entity psi_fix_nch_analog_trigger_tdm is
  generic(ch_nb_g       : natural      := 8;                                              --number of input/output channel
          trig_ext_nb_g : natural      := 1;                                              --number of input external trigger
          fix_fmt_g     : psi_fix_fmt_t:= (1,0,15);                                       --FP format
          rst_pol_g     : std_logic    := '1';                                            -- reset polarity '1' active high
          trig_nb_g     : natural      := 1);                                             --number of output trigger
  port(   clk_i         : in  std_logic;                                                  --processing clock
          rst_i         : in  std_logic;                                                  --Reset  processing '1' <=> active high
          --*** signals ***
          dat_i         : in  std_logic_vector(psi_fix_size(fix_fmt_g)- 1 downto 0);      --// Data Input
          vld_i         : in  std_logic;                                                  --TDM Strobe Input
          ext_i         : in  std_logic_vector(trig_ext_nb_g-1 downto 0);                 --external trigger input
          --*** parameters ***
          mask_min_i    : in std_logic_vector(trig_nb_g*ch_nb_g-1 downto 0);              --mask min results
          mask_max_i    : in std_logic_vector(trig_nb_g*ch_nb_g-1 downto 0);              --mask max results
          mask_ext_i    : in std_logic_vector(trig_nb_g*trig_ext_nb_g-1 downto 0);        --mask external trigger
          thld_min_i    : in std_logic_vector(ch_nb_g*psi_fix_size(fix_fmt_g)-1 downto 0);--thld to set max window
          thld_max_i    : in std_logic_vector(ch_nb_g*psi_fix_size(fix_fmt_g)-1 downto 0);--thld to set Min window
          trig_clr_ext_i: in std_logic_vector(trig_nb_g*trig_ext_nb_g-1 downto 0);
          trig_mode_i   : in std_logic_vector(trig_nb_g-1 downto 0);                      -- Trigger mode (0:Continuous,1:Single) configuration register
          trig_arm_i    : in std_logic_vector(trig_nb_g-1   downto 0);                    -- Arm/dis--arm the trigger, rising edge sensitive
          --*** out ***
          dat_pipe_o    : out std_logic_vector(psi_fix_size(fix_fmt_g)-1 downto 0);       --data out pipelined   for recording
          str_pipe_o    : out std_logic;                                                  --strobe out pipelined for recording
          --*** status ***
          trig_o        : out std_logic_vector(trig_nb_g-1 downto 0);                     --trigger out
          is_arm_o      : out std_logic_vector(trig_nb_g-1 downto 0));                    --trigger is armed
end entity;
--@formatter:on

architecture RTL of psi_fix_nch_analog_trigger_tdm is
  --internal herlpers
  constant len_c          : integer := psi_fix_size(fix_fmt_g);
  type array_thld_t is array (0 to ch_nb_g - 1) of std_logic_vector(len_c - 1 downto 0);
  signal thld_min_array_s : array_thld_t;
  signal thld_max_array_s : array_thld_t;

  type array_mask_t is array (0 to trig_nb_g - 1) of std_logic_vector(ch_nb_g - 1 downto 0);
  signal mask_min_array_s : array_mask_t;
  signal mask_max_array_s : array_mask_t;

  type array_ext_t is array (0 to trig_nb_g - 1) of std_logic_vector(trig_ext_nb_g - 1 downto 0);
  --=================================================================
  -- Comparator mngt signals
  --=================================================================
  signal param_slv2partdm_dat_s : std_logic_vector(ch_nb_g * 2 * len_c - 1 downto 0);
  signal param_slv2partdm_vld_s : std_logic;
  signal str_dff_s              : std_logic;
  signal param_tdm_thld_s       : std_logic_vector(2 * len_c - 1 downto 0);
  signal param_tdm_vld_s        : std_logic;
  signal data_dff0_s            : std_logic_vector(len_c - 1 downto 0);
  signal data_dff1_s            : std_logic_vector(len_c - 1 downto 0);
  signal min_s, max_s, str_s    : std_logic;
  signal min_vector_s           : std_logic_vector(ch_nb_g - 1 downto 0);
  signal max_vector_s           : std_logic_vector(ch_nb_g - 1 downto 0);
  signal comp_str_s             : std_logic;
  --=================================================================
  -- Trigger mngt signals
  --=================================================================
  signal max_trig_s             : array_mask_t; --std_logic_vector(ch_nb_g - 1 downto 0);
  signal min_trig_s             : array_mask_t; --std_logic_vector(ch_nb_g - 1 downto 0);
  signal trig_s                 : std_logic_vector(trig_nb_g - 1 downto 0);
  signal trig_os                : std_logic_vector(trig_nb_g - 1 downto 0);
  --=================================================================
  -- External Trigger mngt signals
  --=================================================================
  signal trig_ext_array_s       : array_ext_t; --external trigger input array
  signal trig_ext_array_dff_s   : array_ext_t; --external trigger input dff array used for edge detect
  signal ext_trig_array_s       : array_ext_t; --external trigger used for trigger
  signal ext_flg_array_s        : array_ext_t; --external trigger flag array
  signal mask_ext_array_s       : array_ext_t;
begin

  --*** helpers construc ***
  gene_mask_trigger_array : for i in 0 to trig_nb_g - 1 generate
  begin
    mask_min_array_s(i) <= mask_min_i((i + 1) * ch_nb_g - 1 downto i * ch_nb_g);
    mask_max_array_s(i) <= mask_max_i((i + 1) * ch_nb_g - 1 downto i * ch_nb_g);
  end generate;

  gene_thld_array : for i in 0 to ch_nb_g - 1 generate
  begin
    thld_min_array_s(i) <= thld_min_i((i + 1) * len_c - 1 downto i * len_c);
    thld_max_array_s(i) <= thld_max_i((i + 1) * len_c - 1 downto i * len_c);
  end generate;

  --*** TAG process dff for input parameter thld ***
  proc_conv_array2slv : process(clk_i)
  begin
    if rising_edge(clk_i) then
      --*** create a big slv to be compatible to further block ***
      for i in 0 to ch_nb_g - 1 loop
        param_slv2partdm_dat_s((i + 1) * 2 * len_c - 1 downto i * 2 * len_c) <= thld_max_array_s(i) & thld_min_array_s(i);
      end loop;
      --*** edge detect ***
      str_dff_s   <= vld_i;
      if vld_i = '1' and str_dff_s = '0' then
        param_slv2partdm_vld_s <= '1';
      else
        param_slv2partdm_vld_s <= '0';
      end if;
      --*** delay 2 stages ***
      data_dff0_s <= dat_i;
      data_dff1_s <= data_dff0_s;
    end if;
  end process;

  --*** TAG inst of parallel to TDM for min/max ***
  inst_par2tdm : entity work.psi_common_par_tdm
    generic map(rst_pol_g  => rst_pol_g,
                ch_nb_g    => ch_nb_g,
                ch_width_g => 2 * len_c)
    port map(                           -- @suppress
      clk_i => clk_i,
      rst_i => rst_i,
      dat_i => param_slv2partdm_dat_s,
      vld_i => param_slv2partdm_vld_s,
      dat_o => param_tdm_thld_s,
      vld_o => param_tdm_vld_s);

  --*** TAG inst of parallel to TDM for min/max ***
  -- 4 stages dff delay
  inst_min_max : entity work.psi_fix_comparator
    generic map(fmt_g     => fix_fmt_g,
                rst_pol_g => rst_pol_g)
    port map(clk_i     => clk_i,
             rst_i     => rst_i,
             set_min_i => param_tdm_thld_s(len_c - 1 downto 0),
             set_max_i => param_tdm_thld_s(2 * len_c - 1 downto len_c),
             data_i    => data_dff1_s,
             vld_i     => param_tdm_vld_s,
             vld_o     => str_s,
             min_o     => min_s,
             max_o     => max_s);

  --*** TAG MASK min with a TDM to parallel for trig gene ***
  inst_tdm_par_min : entity work.psi_common_tdm_par
    generic map(                        
      rst_pol_g => rst_pol_g,
      ch_nb_g => ch_nb_g,
      width_g => 1)
    port map(                           --@suppress
      clk_i    => clk_i,
      rst_i    => rst_i,
      dat_i(0) => min_s,
      vld_i    => str_s,
      dat_o    => min_vector_s,
      vld_o    => open);

  --*** TAG MASK max with a TDM to parallel for trig gene ***
  inst_tdm_par_max : entity work.psi_common_tdm_par
    generic map(                     
      rst_pol_g => rst_pol_g,
      ch_nb_g => ch_nb_g,
      width_g => 1)
    port map(                           --@suppress
      clk_i    => clk_i,
      rst_i    => rst_i,
      dat_i(0) => max_s,
      vld_i    => str_s,
      dat_o    => max_vector_s,
      vld_o    => comp_str_s);

  --*** TAG -> trigger digital from library align data to trigger ***
  inst_delay_data : entity work.psi_common_multi_pl_stage
    generic map(rst_pol_g => rst_pol_g,
                width_g   => len_c,
                use_rdy_g => false,
                stages_g  => 10)
    port map(                           -- @suppress
      clk_i     => clk_i,
      rst_i     => rst_i,
      vld_i     => vld_i,
      dat_i     => dat_i,
      vld_o     => str_pipe_o,
      rdy_i     => '1',
      dat_o     => dat_pipe_o);

  --============================================================================
  -->>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>> TRIGGER MNGT <<<<<<<<<<<<<<<<<<<<<<<<<<<<<
  --============================================================================
  --*** TAG -> MASK **
  proc_mask : process(clk_i)
  begin
    if rising_edge(clk_i) then
      for j in 0 to trig_nb_g - 1 loop
        for i in 0 to ch_nb_g - 1 loop
          if comp_str_s = '1' then
            max_trig_s(j)(i) <= max_vector_s(i) and mask_max_array_s(j)(i);
            min_trig_s(j)(i) <= min_vector_s(i) and mask_min_array_s(j)(i);
          end if;
        end loop;
        -- internal trigger
        if min_trig_s(j) >= to_uslv(1, len_c) or max_trig_s(j) >= to_uslv(1, len_c) or ext_trig_array_s(j) /= to_uslv(0, trig_ext_nb_g) then
          trig_s(j) <= '1';
        else
          trig_s(j) <= '0';
        end if;
      end loop;
    end if;
  end process;

  gene_ext_array : for i in 0 to trig_nb_g - 1 generate
  begin
    trig_ext_array_s(i) <= ext_i;
    mask_ext_array_s(i) <= mask_ext_i((i + 1) * trig_ext_nb_g - 1 downto i * trig_ext_nb_g);
  end generate;

  proc_ext_trig_align : process(clk_i)
  begin
    if rising_edge(clk_i) then
      trig_ext_array_dff_s <= trig_ext_array_s;

      if rst_i = rst_pol_g then
        trig_ext_array_dff_s <= (others => (others => '0'));
        ext_flg_array_s      <= (others => (others => '0'));
      else
        for j in 0 to trig_nb_g - 1 loop
          for k in 0 to trig_ext_nb_g - 1 loop
            --*** rising_edge_detect
            if trig_ext_array_dff_s(j)(k) = '0' and trig_ext_array_s(j)(k) = '1' then
              ext_flg_array_s(j)(k) <= '1';
            elsif trig_clr_ext_i(k) = '1' or trig_os(j) = '1' then
              ext_flg_array_s(j)(k) <= '0';
            end if;
            --*** sync with str
            if comp_str_s = '1' and mask_ext_array_s(j)(k) = '1' then
              ext_trig_array_s(j)(k) <= ext_flg_array_s(j)(k);
            else
              ext_trig_array_s(j)(k) <= '0';
            end if;
          end loop;
        end loop;
      end if;
    end if;
  end process;

  --*** TAG digital trigger from psi common - not the most ressource efficient ***
  gene_trigger_nb : for i in 0 to trig_nb_g - 1 generate
  begin
    inst_trig : entity work.psi_common_trigger_digital
      generic map(trig_nb_g => 1,       --one trigger input
                  rst_pol_g => rst_pol_g) --rst pol set to '1'
      port map(clk_i                       => clk_i, --input clock
               rst_i                       => rst_i, --reset
               trg_mode_cfg_i(0)           => trig_mode_i(i), --single shot mode or continuous
               trg_arm_cfg_i               => trig_arm_i(i), --arming trigger
               trg_edge_cfg_i              => "10", --rising edge forced
               trg_digital_source_cfg_i(0) => '0', --don't care
               digital_trg_i(0)            => trig_s(i), --trigger input
               ext_disarm_i                => '0', --don't care
               trg_is_armed_o              => is_arm_o(i), --trigger status is armed
               trigger_o                   => trig_os(i)); --trigger output
    trig_o <= trig_os;
  end generate;
end architecture;
