------------------------------------------------------------------------------
--  Copyright (c) 2018 by Paul Scherrer Institute, Switzerland
--  All rights reserved.
------------------------------------------------------------------------------

------------------------------------------------------------------------------
-- Libraries
------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
  
library work;
use work.psi_common_array_pkg.all;
  
------------------------------------------------------------------------------
-- Package Declaration
------------------------------------------------------------------------------
package psi_fix_fir_dec_semi_nch_chtdm_conf_rbw_tb_coefs_pkg is

	constant Coefs_R3_48Taps : t_areal(0 to 47) := (
		0.00087738037109375,
		0.001190185546875,
		0.00115203857421875,
		0.00055694580078125,
		-0.00072479248046875,
		-0.0024871826171875,
		-0.003997802734375,
		-0.00415802001953125,
		-0.00202178955078125,
		0.002532958984375,
		0.00824737548828125,
		0.01255035400390625,
		0.0124053955078125,
		0.00576019287109375,
		-0.006988525390625,
		-0.02217864990234375,
		-0.03334808349609375,
		-0.03308868408203125,
		-0.01572418212890625,
		0.020050048828125,
		0.0697784423828125,
		0.12380218505859375,
		0.16971588134765625,
		0.19608306884765625,
		0.19608306884765625,
		0.16971588134765625,
		0.12380218505859375,
		0.0697784423828125,
		0.020050048828125,
		-0.01572418212890625,
		-0.03308868408203125,
		-0.03334808349609375,
		-0.02217864990234375,
		-0.006988525390625,
		0.00576019287109375,
		0.0124053955078125,
		0.01255035400390625,
		0.00824737548828125,
		0.002532958984375,
		-0.00202178955078125,
		-0.00415802001953125,
		-0.003997802734375,
		-0.0024871826171875,
		-0.00072479248046875,
		0.00055694580078125,
		0.00115203857421875,
		0.001190185546875,
		0.00087738037109375);

	constant Coefs_R12_160Taps : t_areal(0 to 159) := (
		-2.288818359375e-05,
		-7.62939453125e-05,
		-0.00012969970703125,
		-0.00018310546875,
		-0.00023651123046875,
		-0.0002899169921875,
		-0.00034332275390625,
		-0.000396728515625,
		-0.0004425048828125,
		-0.00048828125,
		-0.00052642822265625,
		-0.00055694580078125,
		-0.00057220458984375,
		-0.00057220458984375,
		-0.00054931640625,
		-0.00051116943359375,
		-0.0004425048828125,
		-0.0003509521484375,
		-0.0002288818359375,
		-8.392333984375e-05,
		9.1552734375e-05,
		0.0002899169921875,
		0.000518798828125,
		0.000762939453125,
		0.00101470947265625,
		0.00127410888671875,
		0.00153350830078125,
		0.0017852783203125,
		0.00201416015625,
		0.00220489501953125,
		0.00235748291015625,
		0.0024566650390625,
		0.00249481201171875,
		0.00244903564453125,
		0.00232696533203125,
		0.00211334228515625,
		0.00180816650390625,
		0.00141143798828125,
		0.00091552734375,
		0.00032806396484375,
		-0.00034332275390625,
		-0.00109100341796875,
		-0.00189208984375,
		-0.00273895263671875,
		-0.00360107421875,
		-0.00446319580078125,
		-0.00530242919921875,
		-0.00608062744140625,
		-0.00676727294921875,
		-0.00734710693359375,
		-0.007781982421875,
		-0.00803375244140625,
		-0.008087158203125,
		-0.007904052734375,
		-0.007476806640625,
		-0.00677490234375,
		-0.0057830810546875,
		-0.0045013427734375,
		-0.00292205810546875,
		-0.00104522705078125,
		0.0011138916015625,
		0.0035552978515625,
		0.0062408447265625,
		0.0091552734375,
		0.0122528076171875,
		0.0155029296875,
		0.01886749267578125,
		0.0222930908203125,
		0.025726318359375,
		0.02911376953125,
		0.03241729736328125,
		0.0355682373046875,
		0.03852081298828125,
		0.041229248046875,
		0.04364776611328125,
		0.04572296142578125,
		0.04743194580078125,
		0.04874420166015625,
		0.04962921142578125,
		0.05007171630859375,
		0.05007171630859375,
		0.04962921142578125,
		0.04874420166015625,
		0.04743194580078125,
		0.04572296142578125,
		0.04364776611328125,
		0.041229248046875,
		0.03852081298828125,
		0.0355682373046875,
		0.03241729736328125,
		0.02911376953125,
		0.025726318359375,
		0.0222930908203125,
		0.01886749267578125,
		0.0155029296875,
		0.0122528076171875,
		0.0091552734375,
		0.0062408447265625,
		0.0035552978515625,
		0.0011138916015625,
		-0.00104522705078125,
		-0.00292205810546875,
		-0.0045013427734375,
		-0.0057830810546875,
		-0.00677490234375,
		-0.007476806640625,
		-0.007904052734375,
		-0.008087158203125,
		-0.00803375244140625,
		-0.007781982421875,
		-0.00734710693359375,
		-0.00676727294921875,
		-0.00608062744140625,
		-0.00530242919921875,
		-0.00446319580078125,
		-0.00360107421875,
		-0.00273895263671875,
		-0.00189208984375,
		-0.00109100341796875,
		-0.00034332275390625,
		0.00032806396484375,
		0.00091552734375,
		0.00141143798828125,
		0.00180816650390625,
		0.00211334228515625,
		0.00232696533203125,
		0.00244903564453125,
		0.00249481201171875,
		0.0024566650390625,
		0.00235748291015625,
		0.00220489501953125,
		0.00201416015625,
		0.0017852783203125,
		0.00153350830078125,
		0.00127410888671875,
		0.00101470947265625,
		0.000762939453125,
		0.000518798828125,
		0.0002899169921875,
		9.1552734375e-05,
		-8.392333984375e-05,
		-0.0002288818359375,
		-0.0003509521484375,
		-0.0004425048828125,
		-0.00051116943359375,
		-0.00054931640625,
		-0.00057220458984375,
		-0.00057220458984375,
		-0.00055694580078125,
		-0.00052642822265625,
		-0.00048828125,
		-0.0004425048828125,
		-0.000396728515625,
		-0.00034332275390625,
		-0.0002899169921875,
		-0.00023651123046875,
		-0.00018310546875,
		-0.00012969970703125,
		-7.62939453125e-05,
		-2.288818359375e-05);

	constant Coefs_R1_48Taps : t_areal(0 to 47) := (
		0.000335693359375,
		-0.001190185546875,
		0.0004425048828125,
		0.00146484375,
		-0.0019073486328125,
		-0.00095367431640625,
		0.00400543212890625,
		-0.00159454345703125,
		-0.00530242919921875,
		0.00666046142578125,
		0.0031585693359375,
		-0.01258087158203125,
		0.00475311279296875,
		0.01512908935546875,
		-0.018341064453125,
		-0.00849151611328125,
		0.03343963623046875,
		-0.01267242431640625,
		-0.0412750244140625,
		0.0526275634765625,
		0.02672576904296875,
		-0.1241302490234375,
		0.06499481201171875,
		0.51470947265625,
		0.51470947265625,
		0.06499481201171875,
		-0.1241302490234375,
		0.02672576904296875,
		0.0526275634765625,
		-0.0412750244140625,
		-0.01267242431640625,
		0.03343963623046875,
		-0.00849151611328125,
		-0.018341064453125,
		0.01512908935546875,
		0.00475311279296875,
		-0.01258087158203125,
		0.0031585693359375,
		0.00666046142578125,
		-0.00530242919921875,
		-0.00159454345703125,
		0.00400543212890625,
		-0.00095367431640625,
		-0.0019073486328125,
		0.00146484375,
		0.0004425048828125,
		-0.001190185546875,
		0.000335693359375);

end package;

------------------------------------------------------------------------------
-- Package Body
------------------------------------------------------------------------------
package body psi_fix_fir_dec_semi_nch_chtdm_conf_rbw_tb_coefs_pkg is 

end psi_fix_fir_dec_semi_nch_chtdm_conf_rbw_tb_coefs_pkg;
